// soc_system.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        audio_0_external_interface_ADCDAT,                //                  audio_0_external_interface.ADCDAT
		input  wire        audio_0_external_interface_ADCLRCK,               //                                            .ADCLRCK
		input  wire        audio_0_external_interface_BCLK,                  //                                            .BCLK
		output wire        audio_0_external_interface_DACDAT,                //                                            .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,               //                                            .DACLRCK
		inout  wire        audio_and_video_config_0_external_interface_SDAT, // audio_and_video_config_0_external_interface.SDAT
		output wire        audio_and_video_config_0_external_interface_SCLK, //                                            .SCLK
		output wire        audio_pll_0_audio_clk_clk,                        //                       audio_pll_0_audio_clk.clk
		input  wire        clk_clk,                                          //                                         clk.clk
		output wire        hps_hps_io_emac1_inst_TX_CLK,                     //                                         hps.hps_io_emac1_inst_TX_CLK
		output wire        hps_hps_io_emac1_inst_TXD0,                       //                                            .hps_io_emac1_inst_TXD0
		output wire        hps_hps_io_emac1_inst_TXD1,                       //                                            .hps_io_emac1_inst_TXD1
		output wire        hps_hps_io_emac1_inst_TXD2,                       //                                            .hps_io_emac1_inst_TXD2
		output wire        hps_hps_io_emac1_inst_TXD3,                       //                                            .hps_io_emac1_inst_TXD3
		input  wire        hps_hps_io_emac1_inst_RXD0,                       //                                            .hps_io_emac1_inst_RXD0
		inout  wire        hps_hps_io_emac1_inst_MDIO,                       //                                            .hps_io_emac1_inst_MDIO
		output wire        hps_hps_io_emac1_inst_MDC,                        //                                            .hps_io_emac1_inst_MDC
		input  wire        hps_hps_io_emac1_inst_RX_CTL,                     //                                            .hps_io_emac1_inst_RX_CTL
		output wire        hps_hps_io_emac1_inst_TX_CTL,                     //                                            .hps_io_emac1_inst_TX_CTL
		input  wire        hps_hps_io_emac1_inst_RX_CLK,                     //                                            .hps_io_emac1_inst_RX_CLK
		input  wire        hps_hps_io_emac1_inst_RXD1,                       //                                            .hps_io_emac1_inst_RXD1
		input  wire        hps_hps_io_emac1_inst_RXD2,                       //                                            .hps_io_emac1_inst_RXD2
		input  wire        hps_hps_io_emac1_inst_RXD3,                       //                                            .hps_io_emac1_inst_RXD3
		inout  wire        hps_hps_io_sdio_inst_CMD,                         //                                            .hps_io_sdio_inst_CMD
		inout  wire        hps_hps_io_sdio_inst_D0,                          //                                            .hps_io_sdio_inst_D0
		inout  wire        hps_hps_io_sdio_inst_D1,                          //                                            .hps_io_sdio_inst_D1
		output wire        hps_hps_io_sdio_inst_CLK,                         //                                            .hps_io_sdio_inst_CLK
		inout  wire        hps_hps_io_sdio_inst_D2,                          //                                            .hps_io_sdio_inst_D2
		inout  wire        hps_hps_io_sdio_inst_D3,                          //                                            .hps_io_sdio_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D0,                          //                                            .hps_io_usb1_inst_D0
		inout  wire        hps_hps_io_usb1_inst_D1,                          //                                            .hps_io_usb1_inst_D1
		inout  wire        hps_hps_io_usb1_inst_D2,                          //                                            .hps_io_usb1_inst_D2
		inout  wire        hps_hps_io_usb1_inst_D3,                          //                                            .hps_io_usb1_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D4,                          //                                            .hps_io_usb1_inst_D4
		inout  wire        hps_hps_io_usb1_inst_D5,                          //                                            .hps_io_usb1_inst_D5
		inout  wire        hps_hps_io_usb1_inst_D6,                          //                                            .hps_io_usb1_inst_D6
		inout  wire        hps_hps_io_usb1_inst_D7,                          //                                            .hps_io_usb1_inst_D7
		input  wire        hps_hps_io_usb1_inst_CLK,                         //                                            .hps_io_usb1_inst_CLK
		output wire        hps_hps_io_usb1_inst_STP,                         //                                            .hps_io_usb1_inst_STP
		input  wire        hps_hps_io_usb1_inst_DIR,                         //                                            .hps_io_usb1_inst_DIR
		input  wire        hps_hps_io_usb1_inst_NXT,                         //                                            .hps_io_usb1_inst_NXT
		output wire        hps_hps_io_spim1_inst_CLK,                        //                                            .hps_io_spim1_inst_CLK
		output wire        hps_hps_io_spim1_inst_MOSI,                       //                                            .hps_io_spim1_inst_MOSI
		input  wire        hps_hps_io_spim1_inst_MISO,                       //                                            .hps_io_spim1_inst_MISO
		output wire        hps_hps_io_spim1_inst_SS0,                        //                                            .hps_io_spim1_inst_SS0
		input  wire        hps_hps_io_uart0_inst_RX,                         //                                            .hps_io_uart0_inst_RX
		output wire        hps_hps_io_uart0_inst_TX,                         //                                            .hps_io_uart0_inst_TX
		inout  wire        hps_hps_io_i2c0_inst_SDA,                         //                                            .hps_io_i2c0_inst_SDA
		inout  wire        hps_hps_io_i2c0_inst_SCL,                         //                                            .hps_io_i2c0_inst_SCL
		inout  wire        hps_hps_io_i2c1_inst_SDA,                         //                                            .hps_io_i2c1_inst_SDA
		inout  wire        hps_hps_io_i2c1_inst_SCL,                         //                                            .hps_io_i2c1_inst_SCL
		inout  wire        hps_hps_io_gpio_inst_GPIO09,                      //                                            .hps_io_gpio_inst_GPIO09
		inout  wire        hps_hps_io_gpio_inst_GPIO35,                      //                                            .hps_io_gpio_inst_GPIO35
		inout  wire        hps_hps_io_gpio_inst_GPIO40,                      //                                            .hps_io_gpio_inst_GPIO40
		inout  wire        hps_hps_io_gpio_inst_GPIO48,                      //                                            .hps_io_gpio_inst_GPIO48
		inout  wire        hps_hps_io_gpio_inst_GPIO53,                      //                                            .hps_io_gpio_inst_GPIO53
		inout  wire        hps_hps_io_gpio_inst_GPIO54,                      //                                            .hps_io_gpio_inst_GPIO54
		inout  wire        hps_hps_io_gpio_inst_GPIO61,                      //                                            .hps_io_gpio_inst_GPIO61
		output wire [14:0] hps_ddr3_mem_a,                                   //                                    hps_ddr3.mem_a
		output wire [2:0]  hps_ddr3_mem_ba,                                  //                                            .mem_ba
		output wire        hps_ddr3_mem_ck,                                  //                                            .mem_ck
		output wire        hps_ddr3_mem_ck_n,                                //                                            .mem_ck_n
		output wire        hps_ddr3_mem_cke,                                 //                                            .mem_cke
		output wire        hps_ddr3_mem_cs_n,                                //                                            .mem_cs_n
		output wire        hps_ddr3_mem_ras_n,                               //                                            .mem_ras_n
		output wire        hps_ddr3_mem_cas_n,                               //                                            .mem_cas_n
		output wire        hps_ddr3_mem_we_n,                                //                                            .mem_we_n
		output wire        hps_ddr3_mem_reset_n,                             //                                            .mem_reset_n
		inout  wire [31:0] hps_ddr3_mem_dq,                                  //                                            .mem_dq
		inout  wire [3:0]  hps_ddr3_mem_dqs,                                 //                                            .mem_dqs
		inout  wire [3:0]  hps_ddr3_mem_dqs_n,                               //                                            .mem_dqs_n
		output wire        hps_ddr3_mem_odt,                                 //                                            .mem_odt
		output wire [3:0]  hps_ddr3_mem_dm,                                  //                                            .mem_dm
		input  wire        hps_ddr3_oct_rzqin,                               //                                            .oct_rzqin
		input  wire        reset_reset_n,                                    //                                       reset.reset_n
		output wire [7:0]  vga_b,                                            //                                         vga.b
		output wire        vga_blank_n,                                      //                                            .blank_n
		output wire        vga_clk,                                          //                                            .clk
		output wire [7:0]  vga_g,                                            //                                            .g
		output wire        vga_hs,                                           //                                            .hs
		output wire [7:0]  vga_r,                                            //                                            .r
		output wire        vga_sync_n,                                       //                                            .sync_n
		output wire        vga_vs                                            //                                            .vs
	);

	wire         vga_ball_0_avalon_streaming_source_l_valid;             // vga_ball_0:L_VALID -> audio_0:to_dac_left_channel_valid
	wire  [15:0] vga_ball_0_avalon_streaming_source_l_data;              // vga_ball_0:L_DATA -> audio_0:to_dac_left_channel_data
	wire         vga_ball_0_avalon_streaming_source_l_ready;             // audio_0:to_dac_left_channel_ready -> vga_ball_0:L_READY
	wire         vga_ball_0_avalon_streaming_source_r_valid;             // vga_ball_0:R_VALID -> audio_0:to_dac_right_channel_valid
	wire  [15:0] vga_ball_0_avalon_streaming_source_r_data;              // vga_ball_0:R_DATA -> audio_0:to_dac_right_channel_data
	wire         vga_ball_0_avalon_streaming_source_r_ready;             // audio_0:to_dac_right_channel_ready -> vga_ball_0:R_READY
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                        // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                          // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                          // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                         // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                          // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                            // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                        // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                         // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                         // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                         // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                         // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                          // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                        // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                        // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                           // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                         // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                         // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                         // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                        // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                         // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                         // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                          // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                           // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                         // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                        // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_0_vga_ball_0_avalon_slave_0_chipselect; // mm_interconnect_0:vga_ball_0_avalon_slave_0_chipselect -> vga_ball_0:chipselect
	wire   [3:0] mm_interconnect_0_vga_ball_0_avalon_slave_0_address;    // mm_interconnect_0:vga_ball_0_avalon_slave_0_address -> vga_ball_0:address
	wire         mm_interconnect_0_vga_ball_0_avalon_slave_0_write;      // mm_interconnect_0:vga_ball_0_avalon_slave_0_write -> vga_ball_0:write
	wire  [15:0] mm_interconnect_0_vga_ball_0_avalon_slave_0_writedata;  // mm_interconnect_0:vga_ball_0_avalon_slave_0_writedata -> vga_ball_0:writedata
	wire         mm_interconnect_0_p1tank_unit_s1_chipselect;            // mm_interconnect_0:p1tank_unit_s1_chipselect -> p1tank_unit:chipselect
	wire   [7:0] mm_interconnect_0_p1tank_unit_s1_readdata;              // p1tank_unit:readdata -> mm_interconnect_0:p1tank_unit_s1_readdata
	wire         mm_interconnect_0_p1tank_unit_s1_debugaccess;           // mm_interconnect_0:p1tank_unit_s1_debugaccess -> p1tank_unit:debugaccess
	wire  [11:0] mm_interconnect_0_p1tank_unit_s1_address;               // mm_interconnect_0:p1tank_unit_s1_address -> p1tank_unit:address
	wire         mm_interconnect_0_p1tank_unit_s1_write;                 // mm_interconnect_0:p1tank_unit_s1_write -> p1tank_unit:write
	wire   [7:0] mm_interconnect_0_p1tank_unit_s1_writedata;             // mm_interconnect_0:p1tank_unit_s1_writedata -> p1tank_unit:writedata
	wire         mm_interconnect_0_p1tank_unit_s1_clken;                 // mm_interconnect_0:p1tank_unit_s1_clken -> p1tank_unit:clken
	wire         mm_interconnect_0_p2tank_unit_s1_chipselect;            // mm_interconnect_0:p2tank_unit_s1_chipselect -> p2tank_unit:chipselect
	wire   [7:0] mm_interconnect_0_p2tank_unit_s1_readdata;              // p2tank_unit:readdata -> mm_interconnect_0:p2tank_unit_s1_readdata
	wire         mm_interconnect_0_p2tank_unit_s1_debugaccess;           // mm_interconnect_0:p2tank_unit_s1_debugaccess -> p2tank_unit:debugaccess
	wire  [11:0] mm_interconnect_0_p2tank_unit_s1_address;               // mm_interconnect_0:p2tank_unit_s1_address -> p2tank_unit:address
	wire         mm_interconnect_0_p2tank_unit_s1_write;                 // mm_interconnect_0:p2tank_unit_s1_write -> p2tank_unit:write
	wire   [7:0] mm_interconnect_0_p2tank_unit_s1_writedata;             // mm_interconnect_0:p2tank_unit_s1_writedata -> p2tank_unit:writedata
	wire         mm_interconnect_0_p2tank_unit_s1_clken;                 // mm_interconnect_0:p2tank_unit_s1_clken -> p2tank_unit:clken
	wire         mm_interconnect_0_map_unit_s1_chipselect;               // mm_interconnect_0:map_unit_s1_chipselect -> map_unit:chipselect
	wire   [7:0] mm_interconnect_0_map_unit_s1_readdata;                 // map_unit:readdata -> mm_interconnect_0:map_unit_s1_readdata
	wire         mm_interconnect_0_map_unit_s1_debugaccess;              // mm_interconnect_0:map_unit_s1_debugaccess -> map_unit:debugaccess
	wire   [9:0] mm_interconnect_0_map_unit_s1_address;                  // mm_interconnect_0:map_unit_s1_address -> map_unit:address
	wire         mm_interconnect_0_map_unit_s1_write;                    // mm_interconnect_0:map_unit_s1_write -> map_unit:write
	wire   [7:0] mm_interconnect_0_map_unit_s1_writedata;                // mm_interconnect_0:map_unit_s1_writedata -> map_unit:writedata
	wire         mm_interconnect_0_map_unit_s1_clken;                    // mm_interconnect_0:map_unit_s1_clken -> map_unit:clken
	wire         mm_interconnect_0_wall_unit_s1_chipselect;              // mm_interconnect_0:wall_unit_s1_chipselect -> wall_unit:chipselect
	wire   [7:0] mm_interconnect_0_wall_unit_s1_readdata;                // wall_unit:readdata -> mm_interconnect_0:wall_unit_s1_readdata
	wire         mm_interconnect_0_wall_unit_s1_debugaccess;             // mm_interconnect_0:wall_unit_s1_debugaccess -> wall_unit:debugaccess
	wire   [9:0] mm_interconnect_0_wall_unit_s1_address;                 // mm_interconnect_0:wall_unit_s1_address -> wall_unit:address
	wire         mm_interconnect_0_wall_unit_s1_write;                   // mm_interconnect_0:wall_unit_s1_write -> wall_unit:write
	wire   [7:0] mm_interconnect_0_wall_unit_s1_writedata;               // mm_interconnect_0:wall_unit_s1_writedata -> wall_unit:writedata
	wire         mm_interconnect_0_wall_unit_s1_clken;                   // mm_interconnect_0:wall_unit_s1_clken -> wall_unit:clken
	wire         mm_interconnect_0_score_unit_s1_chipselect;             // mm_interconnect_0:score_unit_s1_chipselect -> score_unit:chipselect
	wire   [7:0] mm_interconnect_0_score_unit_s1_readdata;               // score_unit:readdata -> mm_interconnect_0:score_unit_s1_readdata
	wire         mm_interconnect_0_score_unit_s1_debugaccess;            // mm_interconnect_0:score_unit_s1_debugaccess -> score_unit:debugaccess
	wire  [12:0] mm_interconnect_0_score_unit_s1_address;                // mm_interconnect_0:score_unit_s1_address -> score_unit:address
	wire         mm_interconnect_0_score_unit_s1_write;                  // mm_interconnect_0:score_unit_s1_write -> score_unit:write
	wire   [7:0] mm_interconnect_0_score_unit_s1_writedata;              // mm_interconnect_0:score_unit_s1_writedata -> score_unit:writedata
	wire         mm_interconnect_0_score_unit_s1_clken;                  // mm_interconnect_0:score_unit_s1_clken -> score_unit:clken
	wire         mm_interconnect_0_stage_unit_s1_chipselect;             // mm_interconnect_0:stage_unit_s1_chipselect -> stage_unit:chipselect
	wire   [7:0] mm_interconnect_0_stage_unit_s1_readdata;               // stage_unit:readdata -> mm_interconnect_0:stage_unit_s1_readdata
	wire         mm_interconnect_0_stage_unit_s1_debugaccess;            // mm_interconnect_0:stage_unit_s1_debugaccess -> stage_unit:debugaccess
	wire  [10:0] mm_interconnect_0_stage_unit_s1_address;                // mm_interconnect_0:stage_unit_s1_address -> stage_unit:address
	wire         mm_interconnect_0_stage_unit_s1_write;                  // mm_interconnect_0:stage_unit_s1_write -> stage_unit:write
	wire   [7:0] mm_interconnect_0_stage_unit_s1_writedata;              // mm_interconnect_0:stage_unit_s1_writedata -> stage_unit:writedata
	wire         mm_interconnect_0_stage_unit_s1_clken;                  // mm_interconnect_0:stage_unit_s1_clken -> stage_unit:clken
	wire         mm_interconnect_0_num_unit_s1_chipselect;               // mm_interconnect_0:num_unit_s1_chipselect -> num_unit:chipselect
	wire   [7:0] mm_interconnect_0_num_unit_s1_readdata;                 // num_unit:readdata -> mm_interconnect_0:num_unit_s1_readdata
	wire         mm_interconnect_0_num_unit_s1_debugaccess;              // mm_interconnect_0:num_unit_s1_debugaccess -> num_unit:debugaccess
	wire  [10:0] mm_interconnect_0_num_unit_s1_address;                  // mm_interconnect_0:num_unit_s1_address -> num_unit:address
	wire         mm_interconnect_0_num_unit_s1_write;                    // mm_interconnect_0:num_unit_s1_write -> num_unit:write
	wire   [7:0] mm_interconnect_0_num_unit_s1_writedata;                // mm_interconnect_0:num_unit_s1_writedata -> num_unit:writedata
	wire         mm_interconnect_0_num_unit_s1_clken;                    // mm_interconnect_0:num_unit_s1_clken -> num_unit:clken
	wire         mm_interconnect_0_ending_unit_s1_chipselect;            // mm_interconnect_0:ending_unit_s1_chipselect -> ending_unit:chipselect
	wire   [7:0] mm_interconnect_0_ending_unit_s1_readdata;              // ending_unit:readdata -> mm_interconnect_0:ending_unit_s1_readdata
	wire         mm_interconnect_0_ending_unit_s1_debugaccess;           // mm_interconnect_0:ending_unit_s1_debugaccess -> ending_unit:debugaccess
	wire  [10:0] mm_interconnect_0_ending_unit_s1_address;               // mm_interconnect_0:ending_unit_s1_address -> ending_unit:address
	wire         mm_interconnect_0_ending_unit_s1_write;                 // mm_interconnect_0:ending_unit_s1_write -> ending_unit:write
	wire   [7:0] mm_interconnect_0_ending_unit_s1_writedata;             // mm_interconnect_0:ending_unit_s1_writedata -> ending_unit:writedata
	wire         mm_interconnect_0_ending_unit_s1_clken;                 // mm_interconnect_0:ending_unit_s1_clken -> ending_unit:clken
	wire         mm_interconnect_0_explosion_unit_s1_chipselect;         // mm_interconnect_0:explosion_unit_s1_chipselect -> explosion_unit:chipselect
	wire   [7:0] mm_interconnect_0_explosion_unit_s1_readdata;           // explosion_unit:readdata -> mm_interconnect_0:explosion_unit_s1_readdata
	wire         mm_interconnect_0_explosion_unit_s1_debugaccess;        // mm_interconnect_0:explosion_unit_s1_debugaccess -> explosion_unit:debugaccess
	wire  [11:0] mm_interconnect_0_explosion_unit_s1_address;            // mm_interconnect_0:explosion_unit_s1_address -> explosion_unit:address
	wire         mm_interconnect_0_explosion_unit_s1_write;              // mm_interconnect_0:explosion_unit_s1_write -> explosion_unit:write
	wire   [7:0] mm_interconnect_0_explosion_unit_s1_writedata;          // mm_interconnect_0:explosion_unit_s1_writedata -> explosion_unit:writedata
	wire         mm_interconnect_0_explosion_unit_s1_clken;              // mm_interconnect_0:explosion_unit_s1_clken -> explosion_unit:clken
	wire         mm_interconnect_0_jingle_sound_s1_chipselect;           // mm_interconnect_0:jingle_sound_s1_chipselect -> jingle_sound:chipselect
	wire  [15:0] mm_interconnect_0_jingle_sound_s1_readdata;             // jingle_sound:readdata -> mm_interconnect_0:jingle_sound_s1_readdata
	wire         mm_interconnect_0_jingle_sound_s1_debugaccess;          // mm_interconnect_0:jingle_sound_s1_debugaccess -> jingle_sound:debugaccess
	wire  [13:0] mm_interconnect_0_jingle_sound_s1_address;              // mm_interconnect_0:jingle_sound_s1_address -> jingle_sound:address
	wire   [1:0] mm_interconnect_0_jingle_sound_s1_byteenable;           // mm_interconnect_0:jingle_sound_s1_byteenable -> jingle_sound:byteenable
	wire         mm_interconnect_0_jingle_sound_s1_write;                // mm_interconnect_0:jingle_sound_s1_write -> jingle_sound:write
	wire  [15:0] mm_interconnect_0_jingle_sound_s1_writedata;            // mm_interconnect_0:jingle_sound_s1_writedata -> jingle_sound:writedata
	wire         mm_interconnect_0_jingle_sound_s1_clken;                // mm_interconnect_0:jingle_sound_s1_clken -> jingle_sound:clken
	wire         mm_interconnect_0_shoot_sound_s1_chipselect;            // mm_interconnect_0:shoot_sound_s1_chipselect -> shoot_sound:chipselect
	wire  [15:0] mm_interconnect_0_shoot_sound_s1_readdata;              // shoot_sound:readdata -> mm_interconnect_0:shoot_sound_s1_readdata
	wire         mm_interconnect_0_shoot_sound_s1_debugaccess;           // mm_interconnect_0:shoot_sound_s1_debugaccess -> shoot_sound:debugaccess
	wire  [14:0] mm_interconnect_0_shoot_sound_s1_address;               // mm_interconnect_0:shoot_sound_s1_address -> shoot_sound:address
	wire   [1:0] mm_interconnect_0_shoot_sound_s1_byteenable;            // mm_interconnect_0:shoot_sound_s1_byteenable -> shoot_sound:byteenable
	wire         mm_interconnect_0_shoot_sound_s1_write;                 // mm_interconnect_0:shoot_sound_s1_write -> shoot_sound:write
	wire  [15:0] mm_interconnect_0_shoot_sound_s1_writedata;             // mm_interconnect_0:shoot_sound_s1_writedata -> shoot_sound:writedata
	wire         mm_interconnect_0_shoot_sound_s1_clken;                 // mm_interconnect_0:shoot_sound_s1_clken -> shoot_sound:clken
	wire         mm_interconnect_0_crawl_sound_s1_chipselect;            // mm_interconnect_0:crawl_sound_s1_chipselect -> crawl_sound:chipselect
	wire  [15:0] mm_interconnect_0_crawl_sound_s1_readdata;              // crawl_sound:readdata -> mm_interconnect_0:crawl_sound_s1_readdata
	wire         mm_interconnect_0_crawl_sound_s1_debugaccess;           // mm_interconnect_0:crawl_sound_s1_debugaccess -> crawl_sound:debugaccess
	wire  [13:0] mm_interconnect_0_crawl_sound_s1_address;               // mm_interconnect_0:crawl_sound_s1_address -> crawl_sound:address
	wire   [1:0] mm_interconnect_0_crawl_sound_s1_byteenable;            // mm_interconnect_0:crawl_sound_s1_byteenable -> crawl_sound:byteenable
	wire         mm_interconnect_0_crawl_sound_s1_write;                 // mm_interconnect_0:crawl_sound_s1_write -> crawl_sound:write
	wire  [15:0] mm_interconnect_0_crawl_sound_s1_writedata;             // mm_interconnect_0:crawl_sound_s1_writedata -> crawl_sound:writedata
	wire         mm_interconnect_0_crawl_sound_s1_clken;                 // mm_interconnect_0:crawl_sound_s1_clken -> crawl_sound:clken
	wire         mm_interconnect_0_explode_sound_s1_chipselect;          // mm_interconnect_0:explode_sound_s1_chipselect -> explode_sound:chipselect
	wire  [15:0] mm_interconnect_0_explode_sound_s1_readdata;            // explode_sound:readdata -> mm_interconnect_0:explode_sound_s1_readdata
	wire         mm_interconnect_0_explode_sound_s1_debugaccess;         // mm_interconnect_0:explode_sound_s1_debugaccess -> explode_sound:debugaccess
	wire  [13:0] mm_interconnect_0_explode_sound_s1_address;             // mm_interconnect_0:explode_sound_s1_address -> explode_sound:address
	wire   [1:0] mm_interconnect_0_explode_sound_s1_byteenable;          // mm_interconnect_0:explode_sound_s1_byteenable -> explode_sound:byteenable
	wire         mm_interconnect_0_explode_sound_s1_write;               // mm_interconnect_0:explode_sound_s1_write -> explode_sound:write
	wire  [15:0] mm_interconnect_0_explode_sound_s1_writedata;           // mm_interconnect_0:explode_sound_s1_writedata -> explode_sound:writedata
	wire         mm_interconnect_0_explode_sound_s1_clken;               // mm_interconnect_0:explode_sound_s1_clken -> explode_sound:clken
	wire  [31:0] hps_0_f2h_irq0_irq;                                     // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                     // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [audio_0:reset, audio_and_video_config_0:reset, crawl_sound:reset, ending_unit:reset, explode_sound:reset, explosion_unit:reset, jingle_sound:reset, map_unit:reset, mm_interconnect_0:vga_ball_0_reset_reset_bridge_in_reset_reset, num_unit:reset, p1tank_unit:reset, p2tank_unit:reset, rst_translator:in_reset, score_unit:reset, shoot_sound:reset, stage_unit:reset, vga_ball_0:reset, wall_unit:reset]
	wire         rst_controller_reset_out_reset_req;                     // rst_controller:reset_req -> [crawl_sound:reset_req, ending_unit:reset_req, explode_sound:reset_req, explosion_unit:reset_req, jingle_sound:reset_req, map_unit:reset_req, num_unit:reset_req, p1tank_unit:reset_req, p2tank_unit:reset_req, rst_translator:reset_req_in, score_unit:reset_req, shoot_sound:reset_req, stage_unit:reset_req, wall_unit:reset_req]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                                  // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	soc_system_audio_0 audio_0 (
		.clk                          (clk_clk),                                    //                         clk.clk
		.reset                        (rst_controller_reset_out_reset),             //                       reset.reset
		.from_adc_left_channel_ready  (),                                           //  avalon_left_channel_source.ready
		.from_adc_left_channel_data   (),                                           //                            .data
		.from_adc_left_channel_valid  (),                                           //                            .valid
		.from_adc_right_channel_ready (),                                           // avalon_right_channel_source.ready
		.from_adc_right_channel_data  (),                                           //                            .data
		.from_adc_right_channel_valid (),                                           //                            .valid
		.to_dac_left_channel_data     (vga_ball_0_avalon_streaming_source_l_data),  //    avalon_left_channel_sink.data
		.to_dac_left_channel_valid    (vga_ball_0_avalon_streaming_source_l_valid), //                            .valid
		.to_dac_left_channel_ready    (vga_ball_0_avalon_streaming_source_l_ready), //                            .ready
		.to_dac_right_channel_data    (vga_ball_0_avalon_streaming_source_r_data),  //   avalon_right_channel_sink.data
		.to_dac_right_channel_valid   (vga_ball_0_avalon_streaming_source_r_valid), //                            .valid
		.to_dac_right_channel_ready   (vga_ball_0_avalon_streaming_source_r_ready), //                            .ready
		.AUD_ADCDAT                   (audio_0_external_interface_ADCDAT),          //          external_interface.export
		.AUD_ADCLRCK                  (audio_0_external_interface_ADCLRCK),         //                            .export
		.AUD_BCLK                     (audio_0_external_interface_BCLK),            //                            .export
		.AUD_DACDAT                   (audio_0_external_interface_DACDAT),          //                            .export
		.AUD_DACLRCK                  (audio_0_external_interface_DACLRCK)          //                            .export
	);

	soc_system_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clk_clk),                                          //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                   //                  reset.reset
		.address     (),                                                 // avalon_av_config_slave.address
		.byteenable  (),                                                 //                       .byteenable
		.read        (),                                                 //                       .read
		.write       (),                                                 //                       .write
		.writedata   (),                                                 //                       .writedata
		.readdata    (),                                                 //                       .readdata
		.waitrequest (),                                                 //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_0_external_interface_SDAT), //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_0_external_interface_SCLK)  //                       .export
	);

	soc_system_audio_pll_0 audio_pll_0 (
		.ref_clk_clk        (clk_clk),                   //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),            //    ref_reset.reset
		.audio_clk_clk      (audio_pll_0_audio_clk_clk), //    audio_clk.clk
		.reset_source_reset ()                           // reset_source.reset
	);

	soc_system_crawl_sound crawl_sound (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_crawl_sound_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_crawl_sound_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_crawl_sound_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_crawl_sound_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_crawl_sound_s1_write),       //       .write
		.readdata    (mm_interconnect_0_crawl_sound_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_crawl_sound_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_crawl_sound_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	soc_system_ending_unit ending_unit (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_ending_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_ending_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_ending_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_ending_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_ending_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_ending_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_ending_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	soc_system_explode_sound explode_sound (
		.clk         (clk_clk),                                        //   clk1.clk
		.address     (mm_interconnect_0_explode_sound_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_explode_sound_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_explode_sound_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_explode_sound_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_explode_sound_s1_write),       //       .write
		.readdata    (mm_interconnect_0_explode_sound_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_explode_sound_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_explode_sound_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze      (1'b0)                                            // (terminated)
	);

	soc_system_explosion_unit explosion_unit (
		.clk         (clk_clk),                                         //   clk1.clk
		.address     (mm_interconnect_0_explosion_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_explosion_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_explosion_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_explosion_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_explosion_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_explosion_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_explosion_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),                  // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),              //       .reset_req
		.freeze      (1'b0)                                             // (terminated)
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.h2f_user1_clk            (),                                //   h2f_user1_clock.clk
		.mem_a                    (hps_ddr3_mem_a),                  //            memory.mem_a
		.mem_ba                   (hps_ddr3_mem_ba),                 //                  .mem_ba
		.mem_ck                   (hps_ddr3_mem_ck),                 //                  .mem_ck
		.mem_ck_n                 (hps_ddr3_mem_ck_n),               //                  .mem_ck_n
		.mem_cke                  (hps_ddr3_mem_cke),                //                  .mem_cke
		.mem_cs_n                 (hps_ddr3_mem_cs_n),               //                  .mem_cs_n
		.mem_ras_n                (hps_ddr3_mem_ras_n),              //                  .mem_ras_n
		.mem_cas_n                (hps_ddr3_mem_cas_n),              //                  .mem_cas_n
		.mem_we_n                 (hps_ddr3_mem_we_n),               //                  .mem_we_n
		.mem_reset_n              (hps_ddr3_mem_reset_n),            //                  .mem_reset_n
		.mem_dq                   (hps_ddr3_mem_dq),                 //                  .mem_dq
		.mem_dqs                  (hps_ddr3_mem_dqs),                //                  .mem_dqs
		.mem_dqs_n                (hps_ddr3_mem_dqs_n),              //                  .mem_dqs_n
		.mem_odt                  (hps_ddr3_mem_odt),                //                  .mem_odt
		.mem_dm                   (hps_ddr3_mem_dm),                 //                  .mem_dm
		.oct_rzqin                (hps_ddr3_oct_rzqin),              //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_hps_io_emac1_inst_TX_CLK),    //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_hps_io_emac1_inst_TXD0),      //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_hps_io_emac1_inst_TXD1),      //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_hps_io_emac1_inst_TXD2),      //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_hps_io_emac1_inst_TXD3),      //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_hps_io_emac1_inst_RXD0),      //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_hps_io_emac1_inst_MDIO),      //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_hps_io_emac1_inst_MDC),       //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_hps_io_emac1_inst_RX_CTL),    //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_hps_io_emac1_inst_TX_CTL),    //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_hps_io_emac1_inst_RX_CLK),    //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_hps_io_emac1_inst_RXD1),      //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_hps_io_emac1_inst_RXD2),      //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_hps_io_emac1_inst_RXD3),      //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_hps_io_sdio_inst_CMD),        //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_hps_io_sdio_inst_D0),         //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_hps_io_sdio_inst_D1),         //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_hps_io_sdio_inst_CLK),        //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_hps_io_sdio_inst_D2),         //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_hps_io_sdio_inst_D3),         //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_hps_io_usb1_inst_D0),         //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_hps_io_usb1_inst_D1),         //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_hps_io_usb1_inst_D2),         //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_hps_io_usb1_inst_D3),         //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_hps_io_usb1_inst_D4),         //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_hps_io_usb1_inst_D5),         //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_hps_io_usb1_inst_D6),         //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_hps_io_usb1_inst_D7),         //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_hps_io_usb1_inst_CLK),        //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_hps_io_usb1_inst_STP),        //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_hps_io_usb1_inst_DIR),        //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_hps_io_usb1_inst_NXT),        //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_hps_io_spim1_inst_CLK),       //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_hps_io_spim1_inst_MOSI),      //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_hps_io_spim1_inst_MISO),      //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_hps_io_spim1_inst_SS0),       //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_hps_io_uart0_inst_RX),        //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_hps_io_uart0_inst_TX),        //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_hps_io_i2c0_inst_SDA),        //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_hps_io_i2c0_inst_SCL),        //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_hps_io_i2c1_inst_SDA),        //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_hps_io_i2c1_inst_SCL),        //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_hps_io_gpio_inst_GPIO09),     //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_hps_io_gpio_inst_GPIO35),     //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_hps_io_gpio_inst_GPIO40),     //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_hps_io_gpio_inst_GPIO48),     //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_hps_io_gpio_inst_GPIO53),     //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_hps_io_gpio_inst_GPIO54),     //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_hps_io_gpio_inst_GPIO61),     //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                         //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                //                  .awaddr
		.h2f_AWLEN                (),                                //                  .awlen
		.h2f_AWSIZE               (),                                //                  .awsize
		.h2f_AWBURST              (),                                //                  .awburst
		.h2f_AWLOCK               (),                                //                  .awlock
		.h2f_AWCACHE              (),                                //                  .awcache
		.h2f_AWPROT               (),                                //                  .awprot
		.h2f_AWVALID              (),                                //                  .awvalid
		.h2f_AWREADY              (),                                //                  .awready
		.h2f_WID                  (),                                //                  .wid
		.h2f_WDATA                (),                                //                  .wdata
		.h2f_WSTRB                (),                                //                  .wstrb
		.h2f_WLAST                (),                                //                  .wlast
		.h2f_WVALID               (),                                //                  .wvalid
		.h2f_WREADY               (),                                //                  .wready
		.h2f_BID                  (),                                //                  .bid
		.h2f_BRESP                (),                                //                  .bresp
		.h2f_BVALID               (),                                //                  .bvalid
		.h2f_BREADY               (),                                //                  .bready
		.h2f_ARID                 (),                                //                  .arid
		.h2f_ARADDR               (),                                //                  .araddr
		.h2f_ARLEN                (),                                //                  .arlen
		.h2f_ARSIZE               (),                                //                  .arsize
		.h2f_ARBURST              (),                                //                  .arburst
		.h2f_ARLOCK               (),                                //                  .arlock
		.h2f_ARCACHE              (),                                //                  .arcache
		.h2f_ARPROT               (),                                //                  .arprot
		.h2f_ARVALID              (),                                //                  .arvalid
		.h2f_ARREADY              (),                                //                  .arready
		.h2f_RID                  (),                                //                  .rid
		.h2f_RDATA                (),                                //                  .rdata
		.h2f_RRESP                (),                                //                  .rresp
		.h2f_RLAST                (),                                //                  .rlast
		.h2f_RVALID               (),                                //                  .rvalid
		.h2f_RREADY               (),                                //                  .rready
		.f2h_axi_clk              (clk_clk),                         //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                //                  .awaddr
		.f2h_AWLEN                (),                                //                  .awlen
		.f2h_AWSIZE               (),                                //                  .awsize
		.f2h_AWBURST              (),                                //                  .awburst
		.f2h_AWLOCK               (),                                //                  .awlock
		.f2h_AWCACHE              (),                                //                  .awcache
		.f2h_AWPROT               (),                                //                  .awprot
		.f2h_AWVALID              (),                                //                  .awvalid
		.f2h_AWREADY              (),                                //                  .awready
		.f2h_AWUSER               (),                                //                  .awuser
		.f2h_WID                  (),                                //                  .wid
		.f2h_WDATA                (),                                //                  .wdata
		.f2h_WSTRB                (),                                //                  .wstrb
		.f2h_WLAST                (),                                //                  .wlast
		.f2h_WVALID               (),                                //                  .wvalid
		.f2h_WREADY               (),                                //                  .wready
		.f2h_BID                  (),                                //                  .bid
		.f2h_BRESP                (),                                //                  .bresp
		.f2h_BVALID               (),                                //                  .bvalid
		.f2h_BREADY               (),                                //                  .bready
		.f2h_ARID                 (),                                //                  .arid
		.f2h_ARADDR               (),                                //                  .araddr
		.f2h_ARLEN                (),                                //                  .arlen
		.f2h_ARSIZE               (),                                //                  .arsize
		.f2h_ARBURST              (),                                //                  .arburst
		.f2h_ARLOCK               (),                                //                  .arlock
		.f2h_ARCACHE              (),                                //                  .arcache
		.f2h_ARPROT               (),                                //                  .arprot
		.f2h_ARVALID              (),                                //                  .arvalid
		.f2h_ARREADY              (),                                //                  .arready
		.f2h_ARUSER               (),                                //                  .aruser
		.f2h_RID                  (),                                //                  .rid
		.f2h_RDATA                (),                                //                  .rdata
		.f2h_RRESP                (),                                //                  .rresp
		.f2h_RLAST                (),                                //                  .rlast
		.f2h_RVALID               (),                                //                  .rvalid
		.f2h_RREADY               (),                                //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	soc_system_jingle_sound jingle_sound (
		.clk         (clk_clk),                                       //   clk1.clk
		.address     (mm_interconnect_0_jingle_sound_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_jingle_sound_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_jingle_sound_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_jingle_sound_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_jingle_sound_s1_write),       //       .write
		.readdata    (mm_interconnect_0_jingle_sound_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_jingle_sound_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_jingle_sound_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze      (1'b0)                                           // (terminated)
	);

	soc_system_map_unit map_unit (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (mm_interconnect_0_map_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_map_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_map_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_map_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_map_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_map_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_map_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	soc_system_num_unit num_unit (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (mm_interconnect_0_num_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_num_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_num_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_num_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_num_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_num_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_num_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	soc_system_p1tank_unit p1tank_unit (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_p1tank_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p1tank_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p1tank_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p1tank_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p1tank_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p1tank_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p1tank_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	soc_system_p2tank_unit p2tank_unit (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_p2tank_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p2tank_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p2tank_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p2tank_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p2tank_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p2tank_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p2tank_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	soc_system_score_unit score_unit (
		.clk         (clk_clk),                                     //   clk1.clk
		.address     (mm_interconnect_0_score_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_score_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_score_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_score_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_score_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_score_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_score_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	soc_system_shoot_sound shoot_sound (
		.clk         (clk_clk),                                      //   clk1.clk
		.address     (mm_interconnect_0_shoot_sound_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_shoot_sound_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_shoot_sound_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_shoot_sound_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_shoot_sound_s1_write),       //       .write
		.readdata    (mm_interconnect_0_shoot_sound_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_shoot_sound_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_shoot_sound_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),               // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                          // (terminated)
	);

	soc_system_stage_unit stage_unit (
		.clk         (clk_clk),                                     //   clk1.clk
		.address     (mm_interconnect_0_stage_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_stage_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_stage_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_stage_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_stage_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_stage_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_stage_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	vga_ball vga_ball_0 (
		.clk         (clk_clk),                                                //                     clock.clk
		.reset       (rst_controller_reset_out_reset),                         //                     reset.reset
		.writedata   (mm_interconnect_0_vga_ball_0_avalon_slave_0_writedata),  //            avalon_slave_0.writedata
		.write       (mm_interconnect_0_vga_ball_0_avalon_slave_0_write),      //                          .write
		.chipselect  (mm_interconnect_0_vga_ball_0_avalon_slave_0_chipselect), //                          .chipselect
		.address     (mm_interconnect_0_vga_ball_0_avalon_slave_0_address),    //                          .address
		.VGA_B       (vga_b),                                                  //                       vga.b
		.VGA_BLANK_n (vga_blank_n),                                            //                          .blank_n
		.VGA_CLK     (vga_clk),                                                //                          .clk
		.VGA_G       (vga_g),                                                  //                          .g
		.VGA_HS      (vga_hs),                                                 //                          .hs
		.VGA_R       (vga_r),                                                  //                          .r
		.VGA_SYNC_n  (vga_sync_n),                                             //                          .sync_n
		.VGA_VS      (vga_vs),                                                 //                          .vs
		.L_READY     (vga_ball_0_avalon_streaming_source_l_ready),             // avalon_streaming_source_l.ready
		.L_VALID     (vga_ball_0_avalon_streaming_source_l_valid),             //                          .valid
		.L_DATA      (vga_ball_0_avalon_streaming_source_l_data),              //                          .data
		.R_DATA      (vga_ball_0_avalon_streaming_source_r_data),              // avalon_streaming_source_r.data
		.R_READY     (vga_ball_0_avalon_streaming_source_r_ready),             //                          .ready
		.R_VALID     (vga_ball_0_avalon_streaming_source_r_valid)              //                          .valid
	);

	soc_system_wall_unit wall_unit (
		.clk         (clk_clk),                                    //   clk1.clk
		.address     (mm_interconnect_0_wall_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_wall_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_wall_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_wall_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_wall_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_wall_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_wall_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                           //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                         //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                          //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                         //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                        //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                         //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                        //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                         //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                        //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                        //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                            //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                          //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                          //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                          //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                         //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                         //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                            //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                          //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                         //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                         //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                           //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                         //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                          //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                         //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                        //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                         //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                        //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                         //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                        //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                        //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                            //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                          //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                          //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                          //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                         //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                         //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                     // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.vga_ball_0_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                         //                        vga_ball_0_reset_reset_bridge_in_reset.reset
		.crawl_sound_s1_address                                              (mm_interconnect_0_crawl_sound_s1_address),               //                                                crawl_sound_s1.address
		.crawl_sound_s1_write                                                (mm_interconnect_0_crawl_sound_s1_write),                 //                                                              .write
		.crawl_sound_s1_readdata                                             (mm_interconnect_0_crawl_sound_s1_readdata),              //                                                              .readdata
		.crawl_sound_s1_writedata                                            (mm_interconnect_0_crawl_sound_s1_writedata),             //                                                              .writedata
		.crawl_sound_s1_byteenable                                           (mm_interconnect_0_crawl_sound_s1_byteenable),            //                                                              .byteenable
		.crawl_sound_s1_chipselect                                           (mm_interconnect_0_crawl_sound_s1_chipselect),            //                                                              .chipselect
		.crawl_sound_s1_clken                                                (mm_interconnect_0_crawl_sound_s1_clken),                 //                                                              .clken
		.crawl_sound_s1_debugaccess                                          (mm_interconnect_0_crawl_sound_s1_debugaccess),           //                                                              .debugaccess
		.ending_unit_s1_address                                              (mm_interconnect_0_ending_unit_s1_address),               //                                                ending_unit_s1.address
		.ending_unit_s1_write                                                (mm_interconnect_0_ending_unit_s1_write),                 //                                                              .write
		.ending_unit_s1_readdata                                             (mm_interconnect_0_ending_unit_s1_readdata),              //                                                              .readdata
		.ending_unit_s1_writedata                                            (mm_interconnect_0_ending_unit_s1_writedata),             //                                                              .writedata
		.ending_unit_s1_chipselect                                           (mm_interconnect_0_ending_unit_s1_chipselect),            //                                                              .chipselect
		.ending_unit_s1_clken                                                (mm_interconnect_0_ending_unit_s1_clken),                 //                                                              .clken
		.ending_unit_s1_debugaccess                                          (mm_interconnect_0_ending_unit_s1_debugaccess),           //                                                              .debugaccess
		.explode_sound_s1_address                                            (mm_interconnect_0_explode_sound_s1_address),             //                                              explode_sound_s1.address
		.explode_sound_s1_write                                              (mm_interconnect_0_explode_sound_s1_write),               //                                                              .write
		.explode_sound_s1_readdata                                           (mm_interconnect_0_explode_sound_s1_readdata),            //                                                              .readdata
		.explode_sound_s1_writedata                                          (mm_interconnect_0_explode_sound_s1_writedata),           //                                                              .writedata
		.explode_sound_s1_byteenable                                         (mm_interconnect_0_explode_sound_s1_byteenable),          //                                                              .byteenable
		.explode_sound_s1_chipselect                                         (mm_interconnect_0_explode_sound_s1_chipselect),          //                                                              .chipselect
		.explode_sound_s1_clken                                              (mm_interconnect_0_explode_sound_s1_clken),               //                                                              .clken
		.explode_sound_s1_debugaccess                                        (mm_interconnect_0_explode_sound_s1_debugaccess),         //                                                              .debugaccess
		.explosion_unit_s1_address                                           (mm_interconnect_0_explosion_unit_s1_address),            //                                             explosion_unit_s1.address
		.explosion_unit_s1_write                                             (mm_interconnect_0_explosion_unit_s1_write),              //                                                              .write
		.explosion_unit_s1_readdata                                          (mm_interconnect_0_explosion_unit_s1_readdata),           //                                                              .readdata
		.explosion_unit_s1_writedata                                         (mm_interconnect_0_explosion_unit_s1_writedata),          //                                                              .writedata
		.explosion_unit_s1_chipselect                                        (mm_interconnect_0_explosion_unit_s1_chipselect),         //                                                              .chipselect
		.explosion_unit_s1_clken                                             (mm_interconnect_0_explosion_unit_s1_clken),              //                                                              .clken
		.explosion_unit_s1_debugaccess                                       (mm_interconnect_0_explosion_unit_s1_debugaccess),        //                                                              .debugaccess
		.jingle_sound_s1_address                                             (mm_interconnect_0_jingle_sound_s1_address),              //                                               jingle_sound_s1.address
		.jingle_sound_s1_write                                               (mm_interconnect_0_jingle_sound_s1_write),                //                                                              .write
		.jingle_sound_s1_readdata                                            (mm_interconnect_0_jingle_sound_s1_readdata),             //                                                              .readdata
		.jingle_sound_s1_writedata                                           (mm_interconnect_0_jingle_sound_s1_writedata),            //                                                              .writedata
		.jingle_sound_s1_byteenable                                          (mm_interconnect_0_jingle_sound_s1_byteenable),           //                                                              .byteenable
		.jingle_sound_s1_chipselect                                          (mm_interconnect_0_jingle_sound_s1_chipselect),           //                                                              .chipselect
		.jingle_sound_s1_clken                                               (mm_interconnect_0_jingle_sound_s1_clken),                //                                                              .clken
		.jingle_sound_s1_debugaccess                                         (mm_interconnect_0_jingle_sound_s1_debugaccess),          //                                                              .debugaccess
		.map_unit_s1_address                                                 (mm_interconnect_0_map_unit_s1_address),                  //                                                   map_unit_s1.address
		.map_unit_s1_write                                                   (mm_interconnect_0_map_unit_s1_write),                    //                                                              .write
		.map_unit_s1_readdata                                                (mm_interconnect_0_map_unit_s1_readdata),                 //                                                              .readdata
		.map_unit_s1_writedata                                               (mm_interconnect_0_map_unit_s1_writedata),                //                                                              .writedata
		.map_unit_s1_chipselect                                              (mm_interconnect_0_map_unit_s1_chipselect),               //                                                              .chipselect
		.map_unit_s1_clken                                                   (mm_interconnect_0_map_unit_s1_clken),                    //                                                              .clken
		.map_unit_s1_debugaccess                                             (mm_interconnect_0_map_unit_s1_debugaccess),              //                                                              .debugaccess
		.num_unit_s1_address                                                 (mm_interconnect_0_num_unit_s1_address),                  //                                                   num_unit_s1.address
		.num_unit_s1_write                                                   (mm_interconnect_0_num_unit_s1_write),                    //                                                              .write
		.num_unit_s1_readdata                                                (mm_interconnect_0_num_unit_s1_readdata),                 //                                                              .readdata
		.num_unit_s1_writedata                                               (mm_interconnect_0_num_unit_s1_writedata),                //                                                              .writedata
		.num_unit_s1_chipselect                                              (mm_interconnect_0_num_unit_s1_chipselect),               //                                                              .chipselect
		.num_unit_s1_clken                                                   (mm_interconnect_0_num_unit_s1_clken),                    //                                                              .clken
		.num_unit_s1_debugaccess                                             (mm_interconnect_0_num_unit_s1_debugaccess),              //                                                              .debugaccess
		.p1tank_unit_s1_address                                              (mm_interconnect_0_p1tank_unit_s1_address),               //                                                p1tank_unit_s1.address
		.p1tank_unit_s1_write                                                (mm_interconnect_0_p1tank_unit_s1_write),                 //                                                              .write
		.p1tank_unit_s1_readdata                                             (mm_interconnect_0_p1tank_unit_s1_readdata),              //                                                              .readdata
		.p1tank_unit_s1_writedata                                            (mm_interconnect_0_p1tank_unit_s1_writedata),             //                                                              .writedata
		.p1tank_unit_s1_chipselect                                           (mm_interconnect_0_p1tank_unit_s1_chipselect),            //                                                              .chipselect
		.p1tank_unit_s1_clken                                                (mm_interconnect_0_p1tank_unit_s1_clken),                 //                                                              .clken
		.p1tank_unit_s1_debugaccess                                          (mm_interconnect_0_p1tank_unit_s1_debugaccess),           //                                                              .debugaccess
		.p2tank_unit_s1_address                                              (mm_interconnect_0_p2tank_unit_s1_address),               //                                                p2tank_unit_s1.address
		.p2tank_unit_s1_write                                                (mm_interconnect_0_p2tank_unit_s1_write),                 //                                                              .write
		.p2tank_unit_s1_readdata                                             (mm_interconnect_0_p2tank_unit_s1_readdata),              //                                                              .readdata
		.p2tank_unit_s1_writedata                                            (mm_interconnect_0_p2tank_unit_s1_writedata),             //                                                              .writedata
		.p2tank_unit_s1_chipselect                                           (mm_interconnect_0_p2tank_unit_s1_chipselect),            //                                                              .chipselect
		.p2tank_unit_s1_clken                                                (mm_interconnect_0_p2tank_unit_s1_clken),                 //                                                              .clken
		.p2tank_unit_s1_debugaccess                                          (mm_interconnect_0_p2tank_unit_s1_debugaccess),           //                                                              .debugaccess
		.score_unit_s1_address                                               (mm_interconnect_0_score_unit_s1_address),                //                                                 score_unit_s1.address
		.score_unit_s1_write                                                 (mm_interconnect_0_score_unit_s1_write),                  //                                                              .write
		.score_unit_s1_readdata                                              (mm_interconnect_0_score_unit_s1_readdata),               //                                                              .readdata
		.score_unit_s1_writedata                                             (mm_interconnect_0_score_unit_s1_writedata),              //                                                              .writedata
		.score_unit_s1_chipselect                                            (mm_interconnect_0_score_unit_s1_chipselect),             //                                                              .chipselect
		.score_unit_s1_clken                                                 (mm_interconnect_0_score_unit_s1_clken),                  //                                                              .clken
		.score_unit_s1_debugaccess                                           (mm_interconnect_0_score_unit_s1_debugaccess),            //                                                              .debugaccess
		.shoot_sound_s1_address                                              (mm_interconnect_0_shoot_sound_s1_address),               //                                                shoot_sound_s1.address
		.shoot_sound_s1_write                                                (mm_interconnect_0_shoot_sound_s1_write),                 //                                                              .write
		.shoot_sound_s1_readdata                                             (mm_interconnect_0_shoot_sound_s1_readdata),              //                                                              .readdata
		.shoot_sound_s1_writedata                                            (mm_interconnect_0_shoot_sound_s1_writedata),             //                                                              .writedata
		.shoot_sound_s1_byteenable                                           (mm_interconnect_0_shoot_sound_s1_byteenable),            //                                                              .byteenable
		.shoot_sound_s1_chipselect                                           (mm_interconnect_0_shoot_sound_s1_chipselect),            //                                                              .chipselect
		.shoot_sound_s1_clken                                                (mm_interconnect_0_shoot_sound_s1_clken),                 //                                                              .clken
		.shoot_sound_s1_debugaccess                                          (mm_interconnect_0_shoot_sound_s1_debugaccess),           //                                                              .debugaccess
		.stage_unit_s1_address                                               (mm_interconnect_0_stage_unit_s1_address),                //                                                 stage_unit_s1.address
		.stage_unit_s1_write                                                 (mm_interconnect_0_stage_unit_s1_write),                  //                                                              .write
		.stage_unit_s1_readdata                                              (mm_interconnect_0_stage_unit_s1_readdata),               //                                                              .readdata
		.stage_unit_s1_writedata                                             (mm_interconnect_0_stage_unit_s1_writedata),              //                                                              .writedata
		.stage_unit_s1_chipselect                                            (mm_interconnect_0_stage_unit_s1_chipselect),             //                                                              .chipselect
		.stage_unit_s1_clken                                                 (mm_interconnect_0_stage_unit_s1_clken),                  //                                                              .clken
		.stage_unit_s1_debugaccess                                           (mm_interconnect_0_stage_unit_s1_debugaccess),            //                                                              .debugaccess
		.vga_ball_0_avalon_slave_0_address                                   (mm_interconnect_0_vga_ball_0_avalon_slave_0_address),    //                                     vga_ball_0_avalon_slave_0.address
		.vga_ball_0_avalon_slave_0_write                                     (mm_interconnect_0_vga_ball_0_avalon_slave_0_write),      //                                                              .write
		.vga_ball_0_avalon_slave_0_writedata                                 (mm_interconnect_0_vga_ball_0_avalon_slave_0_writedata),  //                                                              .writedata
		.vga_ball_0_avalon_slave_0_chipselect                                (mm_interconnect_0_vga_ball_0_avalon_slave_0_chipselect), //                                                              .chipselect
		.wall_unit_s1_address                                                (mm_interconnect_0_wall_unit_s1_address),                 //                                                  wall_unit_s1.address
		.wall_unit_s1_write                                                  (mm_interconnect_0_wall_unit_s1_write),                   //                                                              .write
		.wall_unit_s1_readdata                                               (mm_interconnect_0_wall_unit_s1_readdata),                //                                                              .readdata
		.wall_unit_s1_writedata                                              (mm_interconnect_0_wall_unit_s1_writedata),               //                                                              .writedata
		.wall_unit_s1_chipselect                                             (mm_interconnect_0_wall_unit_s1_chipselect),              //                                                              .chipselect
		.wall_unit_s1_clken                                                  (mm_interconnect_0_wall_unit_s1_clken),                   //                                                              .clken
		.wall_unit_s1_debugaccess                                            (mm_interconnect_0_wall_unit_s1_debugaccess)              //                                                              .debugaccess
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule

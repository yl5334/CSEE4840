// soc_system.v

// Generated using ACDS version 21.1 842

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        audio_0_external_interface_ADCDAT,                //                  audio_0_external_interface.ADCDAT
		input  wire        audio_0_external_interface_ADCLRCK,               //                                            .ADCLRCK
		input  wire        audio_0_external_interface_BCLK,                  //                                            .BCLK
		output wire        audio_0_external_interface_DACDAT,                //                                            .DACDAT
		input  wire        audio_0_external_interface_DACLRCK,               //                                            .DACLRCK
		inout  wire        audio_and_video_config_0_external_interface_SDAT, // audio_and_video_config_0_external_interface.SDAT
		output wire        audio_and_video_config_0_external_interface_SCLK, //                                            .SCLK
		output wire        audio_pll_0_audio_clk_clk,                        //                       audio_pll_0_audio_clk.clk
		input  wire        clk_clk,                                          //                                         clk.clk
		output wire        hps_hps_io_emac1_inst_TX_CLK,                     //                                         hps.hps_io_emac1_inst_TX_CLK
		output wire        hps_hps_io_emac1_inst_TXD0,                       //                                            .hps_io_emac1_inst_TXD0
		output wire        hps_hps_io_emac1_inst_TXD1,                       //                                            .hps_io_emac1_inst_TXD1
		output wire        hps_hps_io_emac1_inst_TXD2,                       //                                            .hps_io_emac1_inst_TXD2
		output wire        hps_hps_io_emac1_inst_TXD3,                       //                                            .hps_io_emac1_inst_TXD3
		input  wire        hps_hps_io_emac1_inst_RXD0,                       //                                            .hps_io_emac1_inst_RXD0
		inout  wire        hps_hps_io_emac1_inst_MDIO,                       //                                            .hps_io_emac1_inst_MDIO
		output wire        hps_hps_io_emac1_inst_MDC,                        //                                            .hps_io_emac1_inst_MDC
		input  wire        hps_hps_io_emac1_inst_RX_CTL,                     //                                            .hps_io_emac1_inst_RX_CTL
		output wire        hps_hps_io_emac1_inst_TX_CTL,                     //                                            .hps_io_emac1_inst_TX_CTL
		input  wire        hps_hps_io_emac1_inst_RX_CLK,                     //                                            .hps_io_emac1_inst_RX_CLK
		input  wire        hps_hps_io_emac1_inst_RXD1,                       //                                            .hps_io_emac1_inst_RXD1
		input  wire        hps_hps_io_emac1_inst_RXD2,                       //                                            .hps_io_emac1_inst_RXD2
		input  wire        hps_hps_io_emac1_inst_RXD3,                       //                                            .hps_io_emac1_inst_RXD3
		inout  wire        hps_hps_io_sdio_inst_CMD,                         //                                            .hps_io_sdio_inst_CMD
		inout  wire        hps_hps_io_sdio_inst_D0,                          //                                            .hps_io_sdio_inst_D0
		inout  wire        hps_hps_io_sdio_inst_D1,                          //                                            .hps_io_sdio_inst_D1
		output wire        hps_hps_io_sdio_inst_CLK,                         //                                            .hps_io_sdio_inst_CLK
		inout  wire        hps_hps_io_sdio_inst_D2,                          //                                            .hps_io_sdio_inst_D2
		inout  wire        hps_hps_io_sdio_inst_D3,                          //                                            .hps_io_sdio_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D0,                          //                                            .hps_io_usb1_inst_D0
		inout  wire        hps_hps_io_usb1_inst_D1,                          //                                            .hps_io_usb1_inst_D1
		inout  wire        hps_hps_io_usb1_inst_D2,                          //                                            .hps_io_usb1_inst_D2
		inout  wire        hps_hps_io_usb1_inst_D3,                          //                                            .hps_io_usb1_inst_D3
		inout  wire        hps_hps_io_usb1_inst_D4,                          //                                            .hps_io_usb1_inst_D4
		inout  wire        hps_hps_io_usb1_inst_D5,                          //                                            .hps_io_usb1_inst_D5
		inout  wire        hps_hps_io_usb1_inst_D6,                          //                                            .hps_io_usb1_inst_D6
		inout  wire        hps_hps_io_usb1_inst_D7,                          //                                            .hps_io_usb1_inst_D7
		input  wire        hps_hps_io_usb1_inst_CLK,                         //                                            .hps_io_usb1_inst_CLK
		output wire        hps_hps_io_usb1_inst_STP,                         //                                            .hps_io_usb1_inst_STP
		input  wire        hps_hps_io_usb1_inst_DIR,                         //                                            .hps_io_usb1_inst_DIR
		input  wire        hps_hps_io_usb1_inst_NXT,                         //                                            .hps_io_usb1_inst_NXT
		output wire        hps_hps_io_spim1_inst_CLK,                        //                                            .hps_io_spim1_inst_CLK
		output wire        hps_hps_io_spim1_inst_MOSI,                       //                                            .hps_io_spim1_inst_MOSI
		input  wire        hps_hps_io_spim1_inst_MISO,                       //                                            .hps_io_spim1_inst_MISO
		output wire        hps_hps_io_spim1_inst_SS0,                        //                                            .hps_io_spim1_inst_SS0
		input  wire        hps_hps_io_uart0_inst_RX,                         //                                            .hps_io_uart0_inst_RX
		output wire        hps_hps_io_uart0_inst_TX,                         //                                            .hps_io_uart0_inst_TX
		inout  wire        hps_hps_io_i2c0_inst_SDA,                         //                                            .hps_io_i2c0_inst_SDA
		inout  wire        hps_hps_io_i2c0_inst_SCL,                         //                                            .hps_io_i2c0_inst_SCL
		inout  wire        hps_hps_io_i2c1_inst_SDA,                         //                                            .hps_io_i2c1_inst_SDA
		inout  wire        hps_hps_io_i2c1_inst_SCL,                         //                                            .hps_io_i2c1_inst_SCL
		inout  wire        hps_hps_io_gpio_inst_GPIO09,                      //                                            .hps_io_gpio_inst_GPIO09
		inout  wire        hps_hps_io_gpio_inst_GPIO35,                      //                                            .hps_io_gpio_inst_GPIO35
		inout  wire        hps_hps_io_gpio_inst_GPIO40,                      //                                            .hps_io_gpio_inst_GPIO40
		inout  wire        hps_hps_io_gpio_inst_GPIO48,                      //                                            .hps_io_gpio_inst_GPIO48
		inout  wire        hps_hps_io_gpio_inst_GPIO53,                      //                                            .hps_io_gpio_inst_GPIO53
		inout  wire        hps_hps_io_gpio_inst_GPIO54,                      //                                            .hps_io_gpio_inst_GPIO54
		inout  wire        hps_hps_io_gpio_inst_GPIO61,                      //                                            .hps_io_gpio_inst_GPIO61
		output wire [14:0] hps_ddr3_mem_a,                                   //                                    hps_ddr3.mem_a
		output wire [2:0]  hps_ddr3_mem_ba,                                  //                                            .mem_ba
		output wire        hps_ddr3_mem_ck,                                  //                                            .mem_ck
		output wire        hps_ddr3_mem_ck_n,                                //                                            .mem_ck_n
		output wire        hps_ddr3_mem_cke,                                 //                                            .mem_cke
		output wire        hps_ddr3_mem_cs_n,                                //                                            .mem_cs_n
		output wire        hps_ddr3_mem_ras_n,                               //                                            .mem_ras_n
		output wire        hps_ddr3_mem_cas_n,                               //                                            .mem_cas_n
		output wire        hps_ddr3_mem_we_n,                                //                                            .mem_we_n
		output wire        hps_ddr3_mem_reset_n,                             //                                            .mem_reset_n
		inout  wire [31:0] hps_ddr3_mem_dq,                                  //                                            .mem_dq
		inout  wire [3:0]  hps_ddr3_mem_dqs,                                 //                                            .mem_dqs
		inout  wire [3:0]  hps_ddr3_mem_dqs_n,                               //                                            .mem_dqs_n
		output wire        hps_ddr3_mem_odt,                                 //                                            .mem_odt
		output wire [3:0]  hps_ddr3_mem_dm,                                  //                                            .mem_dm
		input  wire        hps_ddr3_oct_rzqin,                               //                                            .oct_rzqin
		input  wire        reset_reset_n,                                    //                                       reset.reset_n
		output wire [7:0]  vga_b,                                            //                                         vga.b
		output wire        vga_blank_n,                                      //                                            .blank_n
		output wire        vga_clk,                                          //                                            .clk
		output wire [7:0]  vga_g,                                            //                                            .g
		output wire        vga_hs,                                           //                                            .hs
		output wire [7:0]  vga_r,                                            //                                            .r
		output wire        vga_sync_n,                                       //                                            .sync_n
		output wire        vga_vs                                            //                                            .vs
	);

	wire         vga_ball_0_avalon_streaming_source_l_valid;             // vga_ball_0:L_VALID -> audio_0:to_dac_left_channel_valid
	wire  [15:0] vga_ball_0_avalon_streaming_source_l_data;              // vga_ball_0:L_DATA -> audio_0:to_dac_left_channel_data
	wire         vga_ball_0_avalon_streaming_source_l_ready;             // audio_0:to_dac_left_channel_ready -> vga_ball_0:L_READY
	wire         vga_ball_0_avalon_streaming_source_r_valid;             // vga_ball_0:R_VALID -> audio_0:to_dac_right_channel_valid
	wire  [15:0] vga_ball_0_avalon_streaming_source_r_data;              // vga_ball_0:R_DATA -> audio_0:to_dac_right_channel_data
	wire         vga_ball_0_avalon_streaming_source_r_ready;             // audio_0:to_dac_right_channel_ready -> vga_ball_0:R_READY
	wire   [1:0] hps_0_h2f_lw_axi_master_awburst;                        // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire   [3:0] hps_0_h2f_lw_axi_master_arlen;                          // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire   [3:0] hps_0_h2f_lw_axi_master_wstrb;                          // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire         hps_0_h2f_lw_axi_master_wready;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire  [11:0] hps_0_h2f_lw_axi_master_rid;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire         hps_0_h2f_lw_axi_master_rready;                         // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire   [3:0] hps_0_h2f_lw_axi_master_awlen;                          // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire  [11:0] hps_0_h2f_lw_axi_master_wid;                            // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire   [3:0] hps_0_h2f_lw_axi_master_arcache;                        // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire         hps_0_h2f_lw_axi_master_wvalid;                         // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_0_h2f_lw_axi_master_araddr;                         // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire   [2:0] hps_0_h2f_lw_axi_master_arprot;                         // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [2:0] hps_0_h2f_lw_axi_master_awprot;                         // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire  [31:0] hps_0_h2f_lw_axi_master_wdata;                          // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire         hps_0_h2f_lw_axi_master_arvalid;                        // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_0_h2f_lw_axi_master_awcache;                        // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire  [11:0] hps_0_h2f_lw_axi_master_arid;                           // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire   [1:0] hps_0_h2f_lw_axi_master_arlock;                         // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire   [1:0] hps_0_h2f_lw_axi_master_awlock;                         // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire  [20:0] hps_0_h2f_lw_axi_master_awaddr;                         // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_0_h2f_lw_axi_master_bresp;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire         hps_0_h2f_lw_axi_master_arready;                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire  [31:0] hps_0_h2f_lw_axi_master_rdata;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire         hps_0_h2f_lw_axi_master_awready;                        // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [1:0] hps_0_h2f_lw_axi_master_arburst;                        // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [2:0] hps_0_h2f_lw_axi_master_arsize;                         // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire         hps_0_h2f_lw_axi_master_bready;                         // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire         hps_0_h2f_lw_axi_master_rlast;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire         hps_0_h2f_lw_axi_master_wlast;                          // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire   [1:0] hps_0_h2f_lw_axi_master_rresp;                          // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire  [11:0] hps_0_h2f_lw_axi_master_awid;                           // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire  [11:0] hps_0_h2f_lw_axi_master_bid;                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire         hps_0_h2f_lw_axi_master_bvalid;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [2:0] hps_0_h2f_lw_axi_master_awsize;                         // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire         hps_0_h2f_lw_axi_master_awvalid;                        // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire         hps_0_h2f_lw_axi_master_rvalid;                         // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire         mm_interconnect_0_vga_ball_0_avalon_slave_0_chipselect; // mm_interconnect_0:vga_ball_0_avalon_slave_0_chipselect -> vga_ball_0:chipselect
	wire   [4:0] mm_interconnect_0_vga_ball_0_avalon_slave_0_address;    // mm_interconnect_0:vga_ball_0_avalon_slave_0_address -> vga_ball_0:address
	wire         mm_interconnect_0_vga_ball_0_avalon_slave_0_write;      // mm_interconnect_0:vga_ball_0_avalon_slave_0_write -> vga_ball_0:write
	wire  [31:0] mm_interconnect_0_vga_ball_0_avalon_slave_0_writedata;  // mm_interconnect_0:vga_ball_0_avalon_slave_0_writedata -> vga_ball_0:writedata
	wire         mm_interconnect_0_p1_unit_s1_chipselect;                // mm_interconnect_0:p1_unit_s1_chipselect -> p1_unit:chipselect
	wire  [15:0] mm_interconnect_0_p1_unit_s1_readdata;                  // p1_unit:readdata -> mm_interconnect_0:p1_unit_s1_readdata
	wire         mm_interconnect_0_p1_unit_s1_debugaccess;               // mm_interconnect_0:p1_unit_s1_debugaccess -> p1_unit:debugaccess
	wire   [9:0] mm_interconnect_0_p1_unit_s1_address;                   // mm_interconnect_0:p1_unit_s1_address -> p1_unit:address
	wire   [1:0] mm_interconnect_0_p1_unit_s1_byteenable;                // mm_interconnect_0:p1_unit_s1_byteenable -> p1_unit:byteenable
	wire         mm_interconnect_0_p1_unit_s1_write;                     // mm_interconnect_0:p1_unit_s1_write -> p1_unit:write
	wire  [15:0] mm_interconnect_0_p1_unit_s1_writedata;                 // mm_interconnect_0:p1_unit_s1_writedata -> p1_unit:writedata
	wire         mm_interconnect_0_p1_unit_s1_clken;                     // mm_interconnect_0:p1_unit_s1_clken -> p1_unit:clken
	wire         mm_interconnect_0_p1_die_s1_chipselect;                 // mm_interconnect_0:p1_die_s1_chipselect -> p1_die:chipselect
	wire  [15:0] mm_interconnect_0_p1_die_s1_readdata;                   // p1_die:readdata -> mm_interconnect_0:p1_die_s1_readdata
	wire         mm_interconnect_0_p1_die_s1_debugaccess;                // mm_interconnect_0:p1_die_s1_debugaccess -> p1_die:debugaccess
	wire   [7:0] mm_interconnect_0_p1_die_s1_address;                    // mm_interconnect_0:p1_die_s1_address -> p1_die:address
	wire   [1:0] mm_interconnect_0_p1_die_s1_byteenable;                 // mm_interconnect_0:p1_die_s1_byteenable -> p1_die:byteenable
	wire         mm_interconnect_0_p1_die_s1_write;                      // mm_interconnect_0:p1_die_s1_write -> p1_die:write
	wire  [15:0] mm_interconnect_0_p1_die_s1_writedata;                  // mm_interconnect_0:p1_die_s1_writedata -> p1_die:writedata
	wire         mm_interconnect_0_p1_die_s1_clken;                      // mm_interconnect_0:p1_die_s1_clken -> p1_die:clken
	wire         mm_interconnect_0_p2_unit_s1_chipselect;                // mm_interconnect_0:p2_unit_s1_chipselect -> p2_unit:chipselect
	wire  [15:0] mm_interconnect_0_p2_unit_s1_readdata;                  // p2_unit:readdata -> mm_interconnect_0:p2_unit_s1_readdata
	wire         mm_interconnect_0_p2_unit_s1_debugaccess;               // mm_interconnect_0:p2_unit_s1_debugaccess -> p2_unit:debugaccess
	wire   [9:0] mm_interconnect_0_p2_unit_s1_address;                   // mm_interconnect_0:p2_unit_s1_address -> p2_unit:address
	wire   [1:0] mm_interconnect_0_p2_unit_s1_byteenable;                // mm_interconnect_0:p2_unit_s1_byteenable -> p2_unit:byteenable
	wire         mm_interconnect_0_p2_unit_s1_write;                     // mm_interconnect_0:p2_unit_s1_write -> p2_unit:write
	wire  [15:0] mm_interconnect_0_p2_unit_s1_writedata;                 // mm_interconnect_0:p2_unit_s1_writedata -> p2_unit:writedata
	wire         mm_interconnect_0_p2_unit_s1_clken;                     // mm_interconnect_0:p2_unit_s1_clken -> p2_unit:clken
	wire         mm_interconnect_0_fix_s1_chipselect;                    // mm_interconnect_0:fix_s1_chipselect -> fix:chipselect
	wire  [15:0] mm_interconnect_0_fix_s1_readdata;                      // fix:readdata -> mm_interconnect_0:fix_s1_readdata
	wire         mm_interconnect_0_fix_s1_debugaccess;                   // mm_interconnect_0:fix_s1_debugaccess -> fix:debugaccess
	wire   [7:0] mm_interconnect_0_fix_s1_address;                       // mm_interconnect_0:fix_s1_address -> fix:address
	wire   [1:0] mm_interconnect_0_fix_s1_byteenable;                    // mm_interconnect_0:fix_s1_byteenable -> fix:byteenable
	wire         mm_interconnect_0_fix_s1_write;                         // mm_interconnect_0:fix_s1_write -> fix:write
	wire  [15:0] mm_interconnect_0_fix_s1_writedata;                     // mm_interconnect_0:fix_s1_writedata -> fix:writedata
	wire         mm_interconnect_0_fix_s1_clken;                         // mm_interconnect_0:fix_s1_clken -> fix:clken
	wire         mm_interconnect_0_bomb_s1_chipselect;                   // mm_interconnect_0:bomb_s1_chipselect -> bomb:chipselect
	wire  [15:0] mm_interconnect_0_bomb_s1_readdata;                     // bomb:readdata -> mm_interconnect_0:bomb_s1_readdata
	wire         mm_interconnect_0_bomb_s1_debugaccess;                  // mm_interconnect_0:bomb_s1_debugaccess -> bomb:debugaccess
	wire   [7:0] mm_interconnect_0_bomb_s1_address;                      // mm_interconnect_0:bomb_s1_address -> bomb:address
	wire   [1:0] mm_interconnect_0_bomb_s1_byteenable;                   // mm_interconnect_0:bomb_s1_byteenable -> bomb:byteenable
	wire         mm_interconnect_0_bomb_s1_write;                        // mm_interconnect_0:bomb_s1_write -> bomb:write
	wire  [15:0] mm_interconnect_0_bomb_s1_writedata;                    // mm_interconnect_0:bomb_s1_writedata -> bomb:writedata
	wire         mm_interconnect_0_bomb_s1_clken;                        // mm_interconnect_0:bomb_s1_clken -> bomb:clken
	wire         mm_interconnect_0_firecenter_s1_chipselect;             // mm_interconnect_0:firecenter_s1_chipselect -> firecenter:chipselect
	wire  [15:0] mm_interconnect_0_firecenter_s1_readdata;               // firecenter:readdata -> mm_interconnect_0:firecenter_s1_readdata
	wire         mm_interconnect_0_firecenter_s1_debugaccess;            // mm_interconnect_0:firecenter_s1_debugaccess -> firecenter:debugaccess
	wire   [7:0] mm_interconnect_0_firecenter_s1_address;                // mm_interconnect_0:firecenter_s1_address -> firecenter:address
	wire   [1:0] mm_interconnect_0_firecenter_s1_byteenable;             // mm_interconnect_0:firecenter_s1_byteenable -> firecenter:byteenable
	wire         mm_interconnect_0_firecenter_s1_write;                  // mm_interconnect_0:firecenter_s1_write -> firecenter:write
	wire  [15:0] mm_interconnect_0_firecenter_s1_writedata;              // mm_interconnect_0:firecenter_s1_writedata -> firecenter:writedata
	wire         mm_interconnect_0_firecenter_s1_clken;                  // mm_interconnect_0:firecenter_s1_clken -> firecenter:clken
	wire         mm_interconnect_0_firehori_s1_chipselect;               // mm_interconnect_0:firehori_s1_chipselect -> firehori:chipselect
	wire  [15:0] mm_interconnect_0_firehori_s1_readdata;                 // firehori:readdata -> mm_interconnect_0:firehori_s1_readdata
	wire         mm_interconnect_0_firehori_s1_debugaccess;              // mm_interconnect_0:firehori_s1_debugaccess -> firehori:debugaccess
	wire   [7:0] mm_interconnect_0_firehori_s1_address;                  // mm_interconnect_0:firehori_s1_address -> firehori:address
	wire   [1:0] mm_interconnect_0_firehori_s1_byteenable;               // mm_interconnect_0:firehori_s1_byteenable -> firehori:byteenable
	wire         mm_interconnect_0_firehori_s1_write;                    // mm_interconnect_0:firehori_s1_write -> firehori:write
	wire  [15:0] mm_interconnect_0_firehori_s1_writedata;                // mm_interconnect_0:firehori_s1_writedata -> firehori:writedata
	wire         mm_interconnect_0_firehori_s1_clken;                    // mm_interconnect_0:firehori_s1_clken -> firehori:clken
	wire         mm_interconnect_0_fireverti_s1_chipselect;              // mm_interconnect_0:fireverti_s1_chipselect -> fireverti:chipselect
	wire  [15:0] mm_interconnect_0_fireverti_s1_readdata;                // fireverti:readdata -> mm_interconnect_0:fireverti_s1_readdata
	wire         mm_interconnect_0_fireverti_s1_debugaccess;             // mm_interconnect_0:fireverti_s1_debugaccess -> fireverti:debugaccess
	wire   [7:0] mm_interconnect_0_fireverti_s1_address;                 // mm_interconnect_0:fireverti_s1_address -> fireverti:address
	wire   [1:0] mm_interconnect_0_fireverti_s1_byteenable;              // mm_interconnect_0:fireverti_s1_byteenable -> fireverti:byteenable
	wire         mm_interconnect_0_fireverti_s1_write;                   // mm_interconnect_0:fireverti_s1_write -> fireverti:write
	wire  [15:0] mm_interconnect_0_fireverti_s1_writedata;               // mm_interconnect_0:fireverti_s1_writedata -> fireverti:writedata
	wire         mm_interconnect_0_fireverti_s1_clken;                   // mm_interconnect_0:fireverti_s1_clken -> fireverti:clken
	wire         mm_interconnect_0_p2_die_s1_chipselect;                 // mm_interconnect_0:p2_die_s1_chipselect -> p2_die:chipselect
	wire  [15:0] mm_interconnect_0_p2_die_s1_readdata;                   // p2_die:readdata -> mm_interconnect_0:p2_die_s1_readdata
	wire         mm_interconnect_0_p2_die_s1_debugaccess;                // mm_interconnect_0:p2_die_s1_debugaccess -> p2_die:debugaccess
	wire   [7:0] mm_interconnect_0_p2_die_s1_address;                    // mm_interconnect_0:p2_die_s1_address -> p2_die:address
	wire   [1:0] mm_interconnect_0_p2_die_s1_byteenable;                 // mm_interconnect_0:p2_die_s1_byteenable -> p2_die:byteenable
	wire         mm_interconnect_0_p2_die_s1_write;                      // mm_interconnect_0:p2_die_s1_write -> p2_die:write
	wire  [15:0] mm_interconnect_0_p2_die_s1_writedata;                  // mm_interconnect_0:p2_die_s1_writedata -> p2_die:writedata
	wire         mm_interconnect_0_p2_die_s1_clken;                      // mm_interconnect_0:p2_die_s1_clken -> p2_die:clken
	wire         mm_interconnect_0_map_unit_s1_chipselect;               // mm_interconnect_0:map_unit_s1_chipselect -> map_unit:chipselect
	wire   [7:0] mm_interconnect_0_map_unit_s1_readdata;                 // map_unit:readdata -> mm_interconnect_0:map_unit_s1_readdata
	wire         mm_interconnect_0_map_unit_s1_debugaccess;              // mm_interconnect_0:map_unit_s1_debugaccess -> map_unit:debugaccess
	wire  [10:0] mm_interconnect_0_map_unit_s1_address;                  // mm_interconnect_0:map_unit_s1_address -> map_unit:address
	wire         mm_interconnect_0_map_unit_s1_write;                    // mm_interconnect_0:map_unit_s1_write -> map_unit:write
	wire   [7:0] mm_interconnect_0_map_unit_s1_writedata;                // mm_interconnect_0:map_unit_s1_writedata -> map_unit:writedata
	wire         mm_interconnect_0_map_unit_s1_clken;                    // mm_interconnect_0:map_unit_s1_clken -> map_unit:clken
	wire         mm_interconnect_0_explode_sound_s1_chipselect;          // mm_interconnect_0:explode_sound_s1_chipselect -> explode_sound:chipselect
	wire  [15:0] mm_interconnect_0_explode_sound_s1_readdata;            // explode_sound:readdata -> mm_interconnect_0:explode_sound_s1_readdata
	wire         mm_interconnect_0_explode_sound_s1_debugaccess;         // mm_interconnect_0:explode_sound_s1_debugaccess -> explode_sound:debugaccess
	wire  [13:0] mm_interconnect_0_explode_sound_s1_address;             // mm_interconnect_0:explode_sound_s1_address -> explode_sound:address
	wire   [1:0] mm_interconnect_0_explode_sound_s1_byteenable;          // mm_interconnect_0:explode_sound_s1_byteenable -> explode_sound:byteenable
	wire         mm_interconnect_0_explode_sound_s1_write;               // mm_interconnect_0:explode_sound_s1_write -> explode_sound:write
	wire  [15:0] mm_interconnect_0_explode_sound_s1_writedata;           // mm_interconnect_0:explode_sound_s1_writedata -> explode_sound:writedata
	wire         mm_interconnect_0_explode_sound_s1_clken;               // mm_interconnect_0:explode_sound_s1_clken -> explode_sound:clken
	wire         mm_interconnect_0_p1_win_s1_chipselect;                 // mm_interconnect_0:p1_win_s1_chipselect -> p1_win:chipselect
	wire  [15:0] mm_interconnect_0_p1_win_s1_readdata;                   // p1_win:readdata -> mm_interconnect_0:p1_win_s1_readdata
	wire         mm_interconnect_0_p1_win_s1_debugaccess;                // mm_interconnect_0:p1_win_s1_debugaccess -> p1_win:debugaccess
	wire  [10:0] mm_interconnect_0_p1_win_s1_address;                    // mm_interconnect_0:p1_win_s1_address -> p1_win:address
	wire   [1:0] mm_interconnect_0_p1_win_s1_byteenable;                 // mm_interconnect_0:p1_win_s1_byteenable -> p1_win:byteenable
	wire         mm_interconnect_0_p1_win_s1_write;                      // mm_interconnect_0:p1_win_s1_write -> p1_win:write
	wire  [15:0] mm_interconnect_0_p1_win_s1_writedata;                  // mm_interconnect_0:p1_win_s1_writedata -> p1_win:writedata
	wire         mm_interconnect_0_p1_win_s1_clken;                      // mm_interconnect_0:p1_win_s1_clken -> p1_win:clken
	wire         mm_interconnect_0_p2_win_s1_chipselect;                 // mm_interconnect_0:p2_win_s1_chipselect -> p2_win:chipselect
	wire  [15:0] mm_interconnect_0_p2_win_s1_readdata;                   // p2_win:readdata -> mm_interconnect_0:p2_win_s1_readdata
	wire         mm_interconnect_0_p2_win_s1_debugaccess;                // mm_interconnect_0:p2_win_s1_debugaccess -> p2_win:debugaccess
	wire  [10:0] mm_interconnect_0_p2_win_s1_address;                    // mm_interconnect_0:p2_win_s1_address -> p2_win:address
	wire   [1:0] mm_interconnect_0_p2_win_s1_byteenable;                 // mm_interconnect_0:p2_win_s1_byteenable -> p2_win:byteenable
	wire         mm_interconnect_0_p2_win_s1_write;                      // mm_interconnect_0:p2_win_s1_write -> p2_win:write
	wire  [15:0] mm_interconnect_0_p2_win_s1_writedata;                  // mm_interconnect_0:p2_win_s1_writedata -> p2_win:writedata
	wire         mm_interconnect_0_p2_win_s1_clken;                      // mm_interconnect_0:p2_win_s1_clken -> p2_win:clken
	wire         mm_interconnect_0_start_s1_chipselect;                  // mm_interconnect_0:start_s1_chipselect -> start:chipselect
	wire  [15:0] mm_interconnect_0_start_s1_readdata;                    // start:readdata -> mm_interconnect_0:start_s1_readdata
	wire         mm_interconnect_0_start_s1_debugaccess;                 // mm_interconnect_0:start_s1_debugaccess -> start:debugaccess
	wire  [11:0] mm_interconnect_0_start_s1_address;                     // mm_interconnect_0:start_s1_address -> start:address
	wire   [1:0] mm_interconnect_0_start_s1_byteenable;                  // mm_interconnect_0:start_s1_byteenable -> start:byteenable
	wire         mm_interconnect_0_start_s1_write;                       // mm_interconnect_0:start_s1_write -> start:write
	wire  [15:0] mm_interconnect_0_start_s1_writedata;                   // mm_interconnect_0:start_s1_writedata -> start:writedata
	wire         mm_interconnect_0_start_s1_clken;                       // mm_interconnect_0:start_s1_clken -> start:clken
	wire         mm_interconnect_0_jingle_sound_s1_chipselect;           // mm_interconnect_0:jingle_sound_s1_chipselect -> jingle_sound:chipselect
	wire  [15:0] mm_interconnect_0_jingle_sound_s1_readdata;             // jingle_sound:readdata -> mm_interconnect_0:jingle_sound_s1_readdata
	wire         mm_interconnect_0_jingle_sound_s1_debugaccess;          // mm_interconnect_0:jingle_sound_s1_debugaccess -> jingle_sound:debugaccess
	wire  [13:0] mm_interconnect_0_jingle_sound_s1_address;              // mm_interconnect_0:jingle_sound_s1_address -> jingle_sound:address
	wire   [1:0] mm_interconnect_0_jingle_sound_s1_byteenable;           // mm_interconnect_0:jingle_sound_s1_byteenable -> jingle_sound:byteenable
	wire         mm_interconnect_0_jingle_sound_s1_write;                // mm_interconnect_0:jingle_sound_s1_write -> jingle_sound:write
	wire  [15:0] mm_interconnect_0_jingle_sound_s1_writedata;            // mm_interconnect_0:jingle_sound_s1_writedata -> jingle_sound:writedata
	wire         mm_interconnect_0_jingle_sound_s1_clken;                // mm_interconnect_0:jingle_sound_s1_clken -> jingle_sound:clken
	wire  [31:0] hps_0_f2h_irq0_irq;                                     // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire  [31:0] hps_0_f2h_irq1_irq;                                     // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire         rst_controller_reset_out_reset;                         // rst_controller:reset_out -> [audio_0:reset, audio_and_video_config_0:reset, bomb:reset, explode_sound:reset, firecenter:reset, firehori:reset, fireverti:reset, fix:reset, jingle_sound:reset, map_unit:reset, mm_interconnect_0:vga_ball_0_reset_reset_bridge_in_reset_reset, p1_die:reset, p1_unit:reset, p1_win:reset, p2_die:reset, p2_unit:reset, p2_win:reset, rst_translator:in_reset, start:reset, vga_ball_0:reset]
	wire         rst_controller_reset_out_reset_req;                     // rst_controller:reset_req -> [bomb:reset_req, explode_sound:reset_req, firecenter:reset_req, firehori:reset_req, fireverti:reset_req, fix:reset_req, jingle_sound:reset_req, map_unit:reset_req, p1_die:reset_req, p1_unit:reset_req, p1_win:reset_req, p2_die:reset_req, p2_unit:reset_req, p2_win:reset_req, rst_translator:reset_req_in, start:reset_req]
	wire         rst_controller_001_reset_out_reset;                     // rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	wire         hps_0_h2f_reset_reset;                                  // hps_0:h2f_rst_n -> rst_controller_001:reset_in0

	soc_system_audio_0 audio_0 (
		.clk                          (clk_clk),                                    //                         clk.clk
		.reset                        (rst_controller_reset_out_reset),             //                       reset.reset
		.from_adc_left_channel_ready  (),                                           //  avalon_left_channel_source.ready
		.from_adc_left_channel_data   (),                                           //                            .data
		.from_adc_left_channel_valid  (),                                           //                            .valid
		.from_adc_right_channel_ready (),                                           // avalon_right_channel_source.ready
		.from_adc_right_channel_data  (),                                           //                            .data
		.from_adc_right_channel_valid (),                                           //                            .valid
		.to_dac_left_channel_data     (vga_ball_0_avalon_streaming_source_l_data),  //    avalon_left_channel_sink.data
		.to_dac_left_channel_valid    (vga_ball_0_avalon_streaming_source_l_valid), //                            .valid
		.to_dac_left_channel_ready    (vga_ball_0_avalon_streaming_source_l_ready), //                            .ready
		.to_dac_right_channel_data    (vga_ball_0_avalon_streaming_source_r_data),  //   avalon_right_channel_sink.data
		.to_dac_right_channel_valid   (vga_ball_0_avalon_streaming_source_r_valid), //                            .valid
		.to_dac_right_channel_ready   (vga_ball_0_avalon_streaming_source_r_ready), //                            .ready
		.AUD_ADCDAT                   (audio_0_external_interface_ADCDAT),          //          external_interface.export
		.AUD_ADCLRCK                  (audio_0_external_interface_ADCLRCK),         //                            .export
		.AUD_BCLK                     (audio_0_external_interface_BCLK),            //                            .export
		.AUD_DACDAT                   (audio_0_external_interface_DACDAT),          //                            .export
		.AUD_DACLRCK                  (audio_0_external_interface_DACLRCK)          //                            .export
	);

	soc_system_audio_and_video_config_0 audio_and_video_config_0 (
		.clk         (clk_clk),                                          //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                   //                  reset.reset
		.address     (),                                                 // avalon_av_config_slave.address
		.byteenable  (),                                                 //                       .byteenable
		.read        (),                                                 //                       .read
		.write       (),                                                 //                       .write
		.writedata   (),                                                 //                       .writedata
		.readdata    (),                                                 //                       .readdata
		.waitrequest (),                                                 //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_0_external_interface_SDAT), //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_0_external_interface_SCLK)  //                       .export
	);

	soc_system_audio_pll_0 audio_pll_0 (
		.ref_clk_clk        (clk_clk),                   //      ref_clk.clk
		.ref_reset_reset    (~reset_reset_n),            //    ref_reset.reset
		.audio_clk_clk      (audio_pll_0_audio_clk_clk), //    audio_clk.clk
		.reset_source_reset ()                           // reset_source.reset
	);

	soc_system_bomb bomb (
		.clk         (clk_clk),                               //   clk1.clk
		.address     (mm_interconnect_0_bomb_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_bomb_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_bomb_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_bomb_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_bomb_s1_write),       //       .write
		.readdata    (mm_interconnect_0_bomb_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_bomb_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_bomb_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),        // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                   // (terminated)
	);

	soc_system_explode_sound explode_sound (
		.clk         (clk_clk),                                        //   clk1.clk
		.address     (mm_interconnect_0_explode_sound_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_explode_sound_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_explode_sound_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_explode_sound_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_explode_sound_s1_write),       //       .write
		.readdata    (mm_interconnect_0_explode_sound_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_explode_sound_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_explode_sound_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze      (1'b0)                                            // (terminated)
	);

	soc_system_firecenter firecenter (
		.clk         (clk_clk),                                     //   clk1.clk
		.address     (mm_interconnect_0_firecenter_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_firecenter_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_firecenter_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_firecenter_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_firecenter_s1_write),       //       .write
		.readdata    (mm_interconnect_0_firecenter_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_firecenter_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_firecenter_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	soc_system_firehori firehori (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (mm_interconnect_0_firehori_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_firehori_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_firehori_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_firehori_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_firehori_s1_write),       //       .write
		.readdata    (mm_interconnect_0_firehori_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_firehori_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_firehori_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	soc_system_fireverti fireverti (
		.clk         (clk_clk),                                    //   clk1.clk
		.address     (mm_interconnect_0_fireverti_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_fireverti_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_fireverti_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_fireverti_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_fireverti_s1_write),       //       .write
		.readdata    (mm_interconnect_0_fireverti_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_fireverti_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_fireverti_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	soc_system_fix fix (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_fix_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_fix_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_fix_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_fix_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_fix_s1_write),       //       .write
		.readdata    (mm_interconnect_0_fix_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_fix_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_fix_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps_0 (
		.h2f_user1_clk            (),                                //   h2f_user1_clock.clk
		.mem_a                    (hps_ddr3_mem_a),                  //            memory.mem_a
		.mem_ba                   (hps_ddr3_mem_ba),                 //                  .mem_ba
		.mem_ck                   (hps_ddr3_mem_ck),                 //                  .mem_ck
		.mem_ck_n                 (hps_ddr3_mem_ck_n),               //                  .mem_ck_n
		.mem_cke                  (hps_ddr3_mem_cke),                //                  .mem_cke
		.mem_cs_n                 (hps_ddr3_mem_cs_n),               //                  .mem_cs_n
		.mem_ras_n                (hps_ddr3_mem_ras_n),              //                  .mem_ras_n
		.mem_cas_n                (hps_ddr3_mem_cas_n),              //                  .mem_cas_n
		.mem_we_n                 (hps_ddr3_mem_we_n),               //                  .mem_we_n
		.mem_reset_n              (hps_ddr3_mem_reset_n),            //                  .mem_reset_n
		.mem_dq                   (hps_ddr3_mem_dq),                 //                  .mem_dq
		.mem_dqs                  (hps_ddr3_mem_dqs),                //                  .mem_dqs
		.mem_dqs_n                (hps_ddr3_mem_dqs_n),              //                  .mem_dqs_n
		.mem_odt                  (hps_ddr3_mem_odt),                //                  .mem_odt
		.mem_dm                   (hps_ddr3_mem_dm),                 //                  .mem_dm
		.oct_rzqin                (hps_ddr3_oct_rzqin),              //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_hps_io_emac1_inst_TX_CLK),    //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_hps_io_emac1_inst_TXD0),      //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_hps_io_emac1_inst_TXD1),      //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_hps_io_emac1_inst_TXD2),      //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_hps_io_emac1_inst_TXD3),      //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_hps_io_emac1_inst_RXD0),      //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_hps_io_emac1_inst_MDIO),      //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_hps_io_emac1_inst_MDC),       //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_hps_io_emac1_inst_RX_CTL),    //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_hps_io_emac1_inst_TX_CTL),    //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_hps_io_emac1_inst_RX_CLK),    //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_hps_io_emac1_inst_RXD1),      //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_hps_io_emac1_inst_RXD2),      //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_hps_io_emac1_inst_RXD3),      //                  .hps_io_emac1_inst_RXD3
		.hps_io_sdio_inst_CMD     (hps_hps_io_sdio_inst_CMD),        //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_hps_io_sdio_inst_D0),         //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_hps_io_sdio_inst_D1),         //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_hps_io_sdio_inst_CLK),        //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_hps_io_sdio_inst_D2),         //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_hps_io_sdio_inst_D3),         //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_hps_io_usb1_inst_D0),         //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_hps_io_usb1_inst_D1),         //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_hps_io_usb1_inst_D2),         //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_hps_io_usb1_inst_D3),         //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_hps_io_usb1_inst_D4),         //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_hps_io_usb1_inst_D5),         //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_hps_io_usb1_inst_D6),         //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_hps_io_usb1_inst_D7),         //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_hps_io_usb1_inst_CLK),        //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_hps_io_usb1_inst_STP),        //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_hps_io_usb1_inst_DIR),        //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_hps_io_usb1_inst_NXT),        //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_hps_io_spim1_inst_CLK),       //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_hps_io_spim1_inst_MOSI),      //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_hps_io_spim1_inst_MISO),      //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_hps_io_spim1_inst_SS0),       //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_hps_io_uart0_inst_RX),        //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_hps_io_uart0_inst_TX),        //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_hps_io_i2c0_inst_SDA),        //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_hps_io_i2c0_inst_SCL),        //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_hps_io_i2c1_inst_SDA),        //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_hps_io_i2c1_inst_SCL),        //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_hps_io_gpio_inst_GPIO09),     //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_hps_io_gpio_inst_GPIO35),     //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_hps_io_gpio_inst_GPIO40),     //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO48  (hps_hps_io_gpio_inst_GPIO48),     //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_hps_io_gpio_inst_GPIO53),     //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_hps_io_gpio_inst_GPIO54),     //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_hps_io_gpio_inst_GPIO61),     //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset),           //         h2f_reset.reset_n
		.h2f_axi_clk              (clk_clk),                         //     h2f_axi_clock.clk
		.h2f_AWID                 (),                                //    h2f_axi_master.awid
		.h2f_AWADDR               (),                                //                  .awaddr
		.h2f_AWLEN                (),                                //                  .awlen
		.h2f_AWSIZE               (),                                //                  .awsize
		.h2f_AWBURST              (),                                //                  .awburst
		.h2f_AWLOCK               (),                                //                  .awlock
		.h2f_AWCACHE              (),                                //                  .awcache
		.h2f_AWPROT               (),                                //                  .awprot
		.h2f_AWVALID              (),                                //                  .awvalid
		.h2f_AWREADY              (),                                //                  .awready
		.h2f_WID                  (),                                //                  .wid
		.h2f_WDATA                (),                                //                  .wdata
		.h2f_WSTRB                (),                                //                  .wstrb
		.h2f_WLAST                (),                                //                  .wlast
		.h2f_WVALID               (),                                //                  .wvalid
		.h2f_WREADY               (),                                //                  .wready
		.h2f_BID                  (),                                //                  .bid
		.h2f_BRESP                (),                                //                  .bresp
		.h2f_BVALID               (),                                //                  .bvalid
		.h2f_BREADY               (),                                //                  .bready
		.h2f_ARID                 (),                                //                  .arid
		.h2f_ARADDR               (),                                //                  .araddr
		.h2f_ARLEN                (),                                //                  .arlen
		.h2f_ARSIZE               (),                                //                  .arsize
		.h2f_ARBURST              (),                                //                  .arburst
		.h2f_ARLOCK               (),                                //                  .arlock
		.h2f_ARCACHE              (),                                //                  .arcache
		.h2f_ARPROT               (),                                //                  .arprot
		.h2f_ARVALID              (),                                //                  .arvalid
		.h2f_ARREADY              (),                                //                  .arready
		.h2f_RID                  (),                                //                  .rid
		.h2f_RDATA                (),                                //                  .rdata
		.h2f_RRESP                (),                                //                  .rresp
		.h2f_RLAST                (),                                //                  .rlast
		.h2f_RVALID               (),                                //                  .rvalid
		.h2f_RREADY               (),                                //                  .rready
		.f2h_axi_clk              (clk_clk),                         //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                //                  .awaddr
		.f2h_AWLEN                (),                                //                  .awlen
		.f2h_AWSIZE               (),                                //                  .awsize
		.f2h_AWBURST              (),                                //                  .awburst
		.f2h_AWLOCK               (),                                //                  .awlock
		.f2h_AWCACHE              (),                                //                  .awcache
		.f2h_AWPROT               (),                                //                  .awprot
		.f2h_AWVALID              (),                                //                  .awvalid
		.f2h_AWREADY              (),                                //                  .awready
		.f2h_AWUSER               (),                                //                  .awuser
		.f2h_WID                  (),                                //                  .wid
		.f2h_WDATA                (),                                //                  .wdata
		.f2h_WSTRB                (),                                //                  .wstrb
		.f2h_WLAST                (),                                //                  .wlast
		.f2h_WVALID               (),                                //                  .wvalid
		.f2h_WREADY               (),                                //                  .wready
		.f2h_BID                  (),                                //                  .bid
		.f2h_BRESP                (),                                //                  .bresp
		.f2h_BVALID               (),                                //                  .bvalid
		.f2h_BREADY               (),                                //                  .bready
		.f2h_ARID                 (),                                //                  .arid
		.f2h_ARADDR               (),                                //                  .araddr
		.f2h_ARLEN                (),                                //                  .arlen
		.f2h_ARSIZE               (),                                //                  .arsize
		.f2h_ARBURST              (),                                //                  .arburst
		.f2h_ARLOCK               (),                                //                  .arlock
		.f2h_ARCACHE              (),                                //                  .arcache
		.f2h_ARPROT               (),                                //                  .arprot
		.f2h_ARVALID              (),                                //                  .arvalid
		.f2h_ARREADY              (),                                //                  .arready
		.f2h_ARUSER               (),                                //                  .aruser
		.f2h_RID                  (),                                //                  .rid
		.f2h_RDATA                (),                                //                  .rdata
		.f2h_RRESP                (),                                //                  .rresp
		.f2h_RLAST                (),                                //                  .rlast
		.f2h_RVALID               (),                                //                  .rvalid
		.f2h_RREADY               (),                                //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                         //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),    // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),  //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),   //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),  //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst), //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),  //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache), //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),  //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid), //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready), //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),     //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),   //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),   //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),   //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),  //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),  //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),     //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),   //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),  //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),  //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),    //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),  //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),   //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),  //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst), //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),  //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache), //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),  //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid), //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready), //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),     //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),   //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),   //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),   //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),  //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),  //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),              //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)               //          f2h_irq1.irq
	);

	soc_system_jingle_sound jingle_sound (
		.clk         (clk_clk),                                       //   clk1.clk
		.address     (mm_interconnect_0_jingle_sound_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_jingle_sound_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_jingle_sound_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_jingle_sound_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_jingle_sound_s1_write),       //       .write
		.readdata    (mm_interconnect_0_jingle_sound_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_jingle_sound_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_jingle_sound_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze      (1'b0)                                           // (terminated)
	);

	soc_system_map_unit map_unit (
		.clk         (clk_clk),                                   //   clk1.clk
		.address     (mm_interconnect_0_map_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_map_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_map_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_map_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_map_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_map_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_map_unit_s1_writedata),   //       .writedata
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	soc_system_p1_die p1_die (
		.clk         (clk_clk),                                 //   clk1.clk
		.address     (mm_interconnect_0_p1_die_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p1_die_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p1_die_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p1_die_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p1_die_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p1_die_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p1_die_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_p1_die_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze      (1'b0)                                     // (terminated)
	);

	soc_system_p1_unit p1_unit (
		.clk         (clk_clk),                                  //   clk1.clk
		.address     (mm_interconnect_0_p1_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p1_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p1_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p1_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p1_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p1_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p1_unit_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_p1_unit_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze      (1'b0)                                      // (terminated)
	);

	soc_system_p1_win p1_win (
		.clk         (clk_clk),                                 //   clk1.clk
		.address     (mm_interconnect_0_p1_win_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p1_win_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p1_win_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p1_win_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p1_win_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p1_win_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p1_win_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_p1_win_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze      (1'b0)                                     // (terminated)
	);

	soc_system_p2_die p2_die (
		.clk         (clk_clk),                                 //   clk1.clk
		.address     (mm_interconnect_0_p2_die_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p2_die_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p2_die_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p2_die_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p2_die_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p2_die_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p2_die_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_p2_die_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze      (1'b0)                                     // (terminated)
	);

	soc_system_p2_unit p2_unit (
		.clk         (clk_clk),                                  //   clk1.clk
		.address     (mm_interconnect_0_p2_unit_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p2_unit_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p2_unit_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p2_unit_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p2_unit_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p2_unit_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p2_unit_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_p2_unit_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),       //       .reset_req
		.freeze      (1'b0)                                      // (terminated)
	);

	soc_system_p2_win p2_win (
		.clk         (clk_clk),                                 //   clk1.clk
		.address     (mm_interconnect_0_p2_win_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_p2_win_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_p2_win_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_p2_win_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_p2_win_s1_write),       //       .write
		.readdata    (mm_interconnect_0_p2_win_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_p2_win_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_p2_win_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),      //       .reset_req
		.freeze      (1'b0)                                     // (terminated)
	);

	soc_system_start start (
		.clk         (clk_clk),                                //   clk1.clk
		.address     (mm_interconnect_0_start_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_start_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_start_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_start_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_start_s1_write),       //       .write
		.readdata    (mm_interconnect_0_start_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_start_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_start_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	vga_ball vga_ball_0 (
		.clk         (clk_clk),                                                //                     clock.clk
		.reset       (rst_controller_reset_out_reset),                         //                     reset.reset
		.writedata   (mm_interconnect_0_vga_ball_0_avalon_slave_0_writedata),  //            avalon_slave_0.writedata
		.write       (mm_interconnect_0_vga_ball_0_avalon_slave_0_write),      //                          .write
		.chipselect  (mm_interconnect_0_vga_ball_0_avalon_slave_0_chipselect), //                          .chipselect
		.address     (mm_interconnect_0_vga_ball_0_avalon_slave_0_address),    //                          .address
		.VGA_B       (vga_b),                                                  //                       vga.b
		.VGA_BLANK_n (vga_blank_n),                                            //                          .blank_n
		.VGA_CLK     (vga_clk),                                                //                          .clk
		.VGA_G       (vga_g),                                                  //                          .g
		.VGA_HS      (vga_hs),                                                 //                          .hs
		.VGA_R       (vga_r),                                                  //                          .r
		.VGA_SYNC_n  (vga_sync_n),                                             //                          .sync_n
		.VGA_VS      (vga_vs),                                                 //                          .vs
		.L_READY     (vga_ball_0_avalon_streaming_source_l_ready),             // avalon_streaming_source_l.ready
		.L_VALID     (vga_ball_0_avalon_streaming_source_l_valid),             //                          .valid
		.L_DATA      (vga_ball_0_avalon_streaming_source_l_data),              //                          .data
		.R_DATA      (vga_ball_0_avalon_streaming_source_r_data),              // avalon_streaming_source_r.data
		.R_READY     (vga_ball_0_avalon_streaming_source_r_ready),             //                          .ready
		.R_VALID     (vga_ball_0_avalon_streaming_source_r_valid)              //                          .valid
	);

	soc_system_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                                        (hps_0_h2f_lw_axi_master_awid),                           //                                       hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                                      (hps_0_h2f_lw_axi_master_awaddr),                         //                                                              .awaddr
		.hps_0_h2f_lw_axi_master_awlen                                       (hps_0_h2f_lw_axi_master_awlen),                          //                                                              .awlen
		.hps_0_h2f_lw_axi_master_awsize                                      (hps_0_h2f_lw_axi_master_awsize),                         //                                                              .awsize
		.hps_0_h2f_lw_axi_master_awburst                                     (hps_0_h2f_lw_axi_master_awburst),                        //                                                              .awburst
		.hps_0_h2f_lw_axi_master_awlock                                      (hps_0_h2f_lw_axi_master_awlock),                         //                                                              .awlock
		.hps_0_h2f_lw_axi_master_awcache                                     (hps_0_h2f_lw_axi_master_awcache),                        //                                                              .awcache
		.hps_0_h2f_lw_axi_master_awprot                                      (hps_0_h2f_lw_axi_master_awprot),                         //                                                              .awprot
		.hps_0_h2f_lw_axi_master_awvalid                                     (hps_0_h2f_lw_axi_master_awvalid),                        //                                                              .awvalid
		.hps_0_h2f_lw_axi_master_awready                                     (hps_0_h2f_lw_axi_master_awready),                        //                                                              .awready
		.hps_0_h2f_lw_axi_master_wid                                         (hps_0_h2f_lw_axi_master_wid),                            //                                                              .wid
		.hps_0_h2f_lw_axi_master_wdata                                       (hps_0_h2f_lw_axi_master_wdata),                          //                                                              .wdata
		.hps_0_h2f_lw_axi_master_wstrb                                       (hps_0_h2f_lw_axi_master_wstrb),                          //                                                              .wstrb
		.hps_0_h2f_lw_axi_master_wlast                                       (hps_0_h2f_lw_axi_master_wlast),                          //                                                              .wlast
		.hps_0_h2f_lw_axi_master_wvalid                                      (hps_0_h2f_lw_axi_master_wvalid),                         //                                                              .wvalid
		.hps_0_h2f_lw_axi_master_wready                                      (hps_0_h2f_lw_axi_master_wready),                         //                                                              .wready
		.hps_0_h2f_lw_axi_master_bid                                         (hps_0_h2f_lw_axi_master_bid),                            //                                                              .bid
		.hps_0_h2f_lw_axi_master_bresp                                       (hps_0_h2f_lw_axi_master_bresp),                          //                                                              .bresp
		.hps_0_h2f_lw_axi_master_bvalid                                      (hps_0_h2f_lw_axi_master_bvalid),                         //                                                              .bvalid
		.hps_0_h2f_lw_axi_master_bready                                      (hps_0_h2f_lw_axi_master_bready),                         //                                                              .bready
		.hps_0_h2f_lw_axi_master_arid                                        (hps_0_h2f_lw_axi_master_arid),                           //                                                              .arid
		.hps_0_h2f_lw_axi_master_araddr                                      (hps_0_h2f_lw_axi_master_araddr),                         //                                                              .araddr
		.hps_0_h2f_lw_axi_master_arlen                                       (hps_0_h2f_lw_axi_master_arlen),                          //                                                              .arlen
		.hps_0_h2f_lw_axi_master_arsize                                      (hps_0_h2f_lw_axi_master_arsize),                         //                                                              .arsize
		.hps_0_h2f_lw_axi_master_arburst                                     (hps_0_h2f_lw_axi_master_arburst),                        //                                                              .arburst
		.hps_0_h2f_lw_axi_master_arlock                                      (hps_0_h2f_lw_axi_master_arlock),                         //                                                              .arlock
		.hps_0_h2f_lw_axi_master_arcache                                     (hps_0_h2f_lw_axi_master_arcache),                        //                                                              .arcache
		.hps_0_h2f_lw_axi_master_arprot                                      (hps_0_h2f_lw_axi_master_arprot),                         //                                                              .arprot
		.hps_0_h2f_lw_axi_master_arvalid                                     (hps_0_h2f_lw_axi_master_arvalid),                        //                                                              .arvalid
		.hps_0_h2f_lw_axi_master_arready                                     (hps_0_h2f_lw_axi_master_arready),                        //                                                              .arready
		.hps_0_h2f_lw_axi_master_rid                                         (hps_0_h2f_lw_axi_master_rid),                            //                                                              .rid
		.hps_0_h2f_lw_axi_master_rdata                                       (hps_0_h2f_lw_axi_master_rdata),                          //                                                              .rdata
		.hps_0_h2f_lw_axi_master_rresp                                       (hps_0_h2f_lw_axi_master_rresp),                          //                                                              .rresp
		.hps_0_h2f_lw_axi_master_rlast                                       (hps_0_h2f_lw_axi_master_rlast),                          //                                                              .rlast
		.hps_0_h2f_lw_axi_master_rvalid                                      (hps_0_h2f_lw_axi_master_rvalid),                         //                                                              .rvalid
		.hps_0_h2f_lw_axi_master_rready                                      (hps_0_h2f_lw_axi_master_rready),                         //                                                              .rready
		.clk_0_clk_clk                                                       (clk_clk),                                                //                                                     clk_0_clk.clk
		.hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                     // hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.vga_ball_0_reset_reset_bridge_in_reset_reset                        (rst_controller_reset_out_reset),                         //                        vga_ball_0_reset_reset_bridge_in_reset.reset
		.bomb_s1_address                                                     (mm_interconnect_0_bomb_s1_address),                      //                                                       bomb_s1.address
		.bomb_s1_write                                                       (mm_interconnect_0_bomb_s1_write),                        //                                                              .write
		.bomb_s1_readdata                                                    (mm_interconnect_0_bomb_s1_readdata),                     //                                                              .readdata
		.bomb_s1_writedata                                                   (mm_interconnect_0_bomb_s1_writedata),                    //                                                              .writedata
		.bomb_s1_byteenable                                                  (mm_interconnect_0_bomb_s1_byteenable),                   //                                                              .byteenable
		.bomb_s1_chipselect                                                  (mm_interconnect_0_bomb_s1_chipselect),                   //                                                              .chipselect
		.bomb_s1_clken                                                       (mm_interconnect_0_bomb_s1_clken),                        //                                                              .clken
		.bomb_s1_debugaccess                                                 (mm_interconnect_0_bomb_s1_debugaccess),                  //                                                              .debugaccess
		.explode_sound_s1_address                                            (mm_interconnect_0_explode_sound_s1_address),             //                                              explode_sound_s1.address
		.explode_sound_s1_write                                              (mm_interconnect_0_explode_sound_s1_write),               //                                                              .write
		.explode_sound_s1_readdata                                           (mm_interconnect_0_explode_sound_s1_readdata),            //                                                              .readdata
		.explode_sound_s1_writedata                                          (mm_interconnect_0_explode_sound_s1_writedata),           //                                                              .writedata
		.explode_sound_s1_byteenable                                         (mm_interconnect_0_explode_sound_s1_byteenable),          //                                                              .byteenable
		.explode_sound_s1_chipselect                                         (mm_interconnect_0_explode_sound_s1_chipselect),          //                                                              .chipselect
		.explode_sound_s1_clken                                              (mm_interconnect_0_explode_sound_s1_clken),               //                                                              .clken
		.explode_sound_s1_debugaccess                                        (mm_interconnect_0_explode_sound_s1_debugaccess),         //                                                              .debugaccess
		.firecenter_s1_address                                               (mm_interconnect_0_firecenter_s1_address),                //                                                 firecenter_s1.address
		.firecenter_s1_write                                                 (mm_interconnect_0_firecenter_s1_write),                  //                                                              .write
		.firecenter_s1_readdata                                              (mm_interconnect_0_firecenter_s1_readdata),               //                                                              .readdata
		.firecenter_s1_writedata                                             (mm_interconnect_0_firecenter_s1_writedata),              //                                                              .writedata
		.firecenter_s1_byteenable                                            (mm_interconnect_0_firecenter_s1_byteenable),             //                                                              .byteenable
		.firecenter_s1_chipselect                                            (mm_interconnect_0_firecenter_s1_chipselect),             //                                                              .chipselect
		.firecenter_s1_clken                                                 (mm_interconnect_0_firecenter_s1_clken),                  //                                                              .clken
		.firecenter_s1_debugaccess                                           (mm_interconnect_0_firecenter_s1_debugaccess),            //                                                              .debugaccess
		.firehori_s1_address                                                 (mm_interconnect_0_firehori_s1_address),                  //                                                   firehori_s1.address
		.firehori_s1_write                                                   (mm_interconnect_0_firehori_s1_write),                    //                                                              .write
		.firehori_s1_readdata                                                (mm_interconnect_0_firehori_s1_readdata),                 //                                                              .readdata
		.firehori_s1_writedata                                               (mm_interconnect_0_firehori_s1_writedata),                //                                                              .writedata
		.firehori_s1_byteenable                                              (mm_interconnect_0_firehori_s1_byteenable),               //                                                              .byteenable
		.firehori_s1_chipselect                                              (mm_interconnect_0_firehori_s1_chipselect),               //                                                              .chipselect
		.firehori_s1_clken                                                   (mm_interconnect_0_firehori_s1_clken),                    //                                                              .clken
		.firehori_s1_debugaccess                                             (mm_interconnect_0_firehori_s1_debugaccess),              //                                                              .debugaccess
		.fireverti_s1_address                                                (mm_interconnect_0_fireverti_s1_address),                 //                                                  fireverti_s1.address
		.fireverti_s1_write                                                  (mm_interconnect_0_fireverti_s1_write),                   //                                                              .write
		.fireverti_s1_readdata                                               (mm_interconnect_0_fireverti_s1_readdata),                //                                                              .readdata
		.fireverti_s1_writedata                                              (mm_interconnect_0_fireverti_s1_writedata),               //                                                              .writedata
		.fireverti_s1_byteenable                                             (mm_interconnect_0_fireverti_s1_byteenable),              //                                                              .byteenable
		.fireverti_s1_chipselect                                             (mm_interconnect_0_fireverti_s1_chipselect),              //                                                              .chipselect
		.fireverti_s1_clken                                                  (mm_interconnect_0_fireverti_s1_clken),                   //                                                              .clken
		.fireverti_s1_debugaccess                                            (mm_interconnect_0_fireverti_s1_debugaccess),             //                                                              .debugaccess
		.fix_s1_address                                                      (mm_interconnect_0_fix_s1_address),                       //                                                        fix_s1.address
		.fix_s1_write                                                        (mm_interconnect_0_fix_s1_write),                         //                                                              .write
		.fix_s1_readdata                                                     (mm_interconnect_0_fix_s1_readdata),                      //                                                              .readdata
		.fix_s1_writedata                                                    (mm_interconnect_0_fix_s1_writedata),                     //                                                              .writedata
		.fix_s1_byteenable                                                   (mm_interconnect_0_fix_s1_byteenable),                    //                                                              .byteenable
		.fix_s1_chipselect                                                   (mm_interconnect_0_fix_s1_chipselect),                    //                                                              .chipselect
		.fix_s1_clken                                                        (mm_interconnect_0_fix_s1_clken),                         //                                                              .clken
		.fix_s1_debugaccess                                                  (mm_interconnect_0_fix_s1_debugaccess),                   //                                                              .debugaccess
		.jingle_sound_s1_address                                             (mm_interconnect_0_jingle_sound_s1_address),              //                                               jingle_sound_s1.address
		.jingle_sound_s1_write                                               (mm_interconnect_0_jingle_sound_s1_write),                //                                                              .write
		.jingle_sound_s1_readdata                                            (mm_interconnect_0_jingle_sound_s1_readdata),             //                                                              .readdata
		.jingle_sound_s1_writedata                                           (mm_interconnect_0_jingle_sound_s1_writedata),            //                                                              .writedata
		.jingle_sound_s1_byteenable                                          (mm_interconnect_0_jingle_sound_s1_byteenable),           //                                                              .byteenable
		.jingle_sound_s1_chipselect                                          (mm_interconnect_0_jingle_sound_s1_chipselect),           //                                                              .chipselect
		.jingle_sound_s1_clken                                               (mm_interconnect_0_jingle_sound_s1_clken),                //                                                              .clken
		.jingle_sound_s1_debugaccess                                         (mm_interconnect_0_jingle_sound_s1_debugaccess),          //                                                              .debugaccess
		.map_unit_s1_address                                                 (mm_interconnect_0_map_unit_s1_address),                  //                                                   map_unit_s1.address
		.map_unit_s1_write                                                   (mm_interconnect_0_map_unit_s1_write),                    //                                                              .write
		.map_unit_s1_readdata                                                (mm_interconnect_0_map_unit_s1_readdata),                 //                                                              .readdata
		.map_unit_s1_writedata                                               (mm_interconnect_0_map_unit_s1_writedata),                //                                                              .writedata
		.map_unit_s1_chipselect                                              (mm_interconnect_0_map_unit_s1_chipselect),               //                                                              .chipselect
		.map_unit_s1_clken                                                   (mm_interconnect_0_map_unit_s1_clken),                    //                                                              .clken
		.map_unit_s1_debugaccess                                             (mm_interconnect_0_map_unit_s1_debugaccess),              //                                                              .debugaccess
		.p1_die_s1_address                                                   (mm_interconnect_0_p1_die_s1_address),                    //                                                     p1_die_s1.address
		.p1_die_s1_write                                                     (mm_interconnect_0_p1_die_s1_write),                      //                                                              .write
		.p1_die_s1_readdata                                                  (mm_interconnect_0_p1_die_s1_readdata),                   //                                                              .readdata
		.p1_die_s1_writedata                                                 (mm_interconnect_0_p1_die_s1_writedata),                  //                                                              .writedata
		.p1_die_s1_byteenable                                                (mm_interconnect_0_p1_die_s1_byteenable),                 //                                                              .byteenable
		.p1_die_s1_chipselect                                                (mm_interconnect_0_p1_die_s1_chipselect),                 //                                                              .chipselect
		.p1_die_s1_clken                                                     (mm_interconnect_0_p1_die_s1_clken),                      //                                                              .clken
		.p1_die_s1_debugaccess                                               (mm_interconnect_0_p1_die_s1_debugaccess),                //                                                              .debugaccess
		.p1_unit_s1_address                                                  (mm_interconnect_0_p1_unit_s1_address),                   //                                                    p1_unit_s1.address
		.p1_unit_s1_write                                                    (mm_interconnect_0_p1_unit_s1_write),                     //                                                              .write
		.p1_unit_s1_readdata                                                 (mm_interconnect_0_p1_unit_s1_readdata),                  //                                                              .readdata
		.p1_unit_s1_writedata                                                (mm_interconnect_0_p1_unit_s1_writedata),                 //                                                              .writedata
		.p1_unit_s1_byteenable                                               (mm_interconnect_0_p1_unit_s1_byteenable),                //                                                              .byteenable
		.p1_unit_s1_chipselect                                               (mm_interconnect_0_p1_unit_s1_chipselect),                //                                                              .chipselect
		.p1_unit_s1_clken                                                    (mm_interconnect_0_p1_unit_s1_clken),                     //                                                              .clken
		.p1_unit_s1_debugaccess                                              (mm_interconnect_0_p1_unit_s1_debugaccess),               //                                                              .debugaccess
		.p1_win_s1_address                                                   (mm_interconnect_0_p1_win_s1_address),                    //                                                     p1_win_s1.address
		.p1_win_s1_write                                                     (mm_interconnect_0_p1_win_s1_write),                      //                                                              .write
		.p1_win_s1_readdata                                                  (mm_interconnect_0_p1_win_s1_readdata),                   //                                                              .readdata
		.p1_win_s1_writedata                                                 (mm_interconnect_0_p1_win_s1_writedata),                  //                                                              .writedata
		.p1_win_s1_byteenable                                                (mm_interconnect_0_p1_win_s1_byteenable),                 //                                                              .byteenable
		.p1_win_s1_chipselect                                                (mm_interconnect_0_p1_win_s1_chipselect),                 //                                                              .chipselect
		.p1_win_s1_clken                                                     (mm_interconnect_0_p1_win_s1_clken),                      //                                                              .clken
		.p1_win_s1_debugaccess                                               (mm_interconnect_0_p1_win_s1_debugaccess),                //                                                              .debugaccess
		.p2_die_s1_address                                                   (mm_interconnect_0_p2_die_s1_address),                    //                                                     p2_die_s1.address
		.p2_die_s1_write                                                     (mm_interconnect_0_p2_die_s1_write),                      //                                                              .write
		.p2_die_s1_readdata                                                  (mm_interconnect_0_p2_die_s1_readdata),                   //                                                              .readdata
		.p2_die_s1_writedata                                                 (mm_interconnect_0_p2_die_s1_writedata),                  //                                                              .writedata
		.p2_die_s1_byteenable                                                (mm_interconnect_0_p2_die_s1_byteenable),                 //                                                              .byteenable
		.p2_die_s1_chipselect                                                (mm_interconnect_0_p2_die_s1_chipselect),                 //                                                              .chipselect
		.p2_die_s1_clken                                                     (mm_interconnect_0_p2_die_s1_clken),                      //                                                              .clken
		.p2_die_s1_debugaccess                                               (mm_interconnect_0_p2_die_s1_debugaccess),                //                                                              .debugaccess
		.p2_unit_s1_address                                                  (mm_interconnect_0_p2_unit_s1_address),                   //                                                    p2_unit_s1.address
		.p2_unit_s1_write                                                    (mm_interconnect_0_p2_unit_s1_write),                     //                                                              .write
		.p2_unit_s1_readdata                                                 (mm_interconnect_0_p2_unit_s1_readdata),                  //                                                              .readdata
		.p2_unit_s1_writedata                                                (mm_interconnect_0_p2_unit_s1_writedata),                 //                                                              .writedata
		.p2_unit_s1_byteenable                                               (mm_interconnect_0_p2_unit_s1_byteenable),                //                                                              .byteenable
		.p2_unit_s1_chipselect                                               (mm_interconnect_0_p2_unit_s1_chipselect),                //                                                              .chipselect
		.p2_unit_s1_clken                                                    (mm_interconnect_0_p2_unit_s1_clken),                     //                                                              .clken
		.p2_unit_s1_debugaccess                                              (mm_interconnect_0_p2_unit_s1_debugaccess),               //                                                              .debugaccess
		.p2_win_s1_address                                                   (mm_interconnect_0_p2_win_s1_address),                    //                                                     p2_win_s1.address
		.p2_win_s1_write                                                     (mm_interconnect_0_p2_win_s1_write),                      //                                                              .write
		.p2_win_s1_readdata                                                  (mm_interconnect_0_p2_win_s1_readdata),                   //                                                              .readdata
		.p2_win_s1_writedata                                                 (mm_interconnect_0_p2_win_s1_writedata),                  //                                                              .writedata
		.p2_win_s1_byteenable                                                (mm_interconnect_0_p2_win_s1_byteenable),                 //                                                              .byteenable
		.p2_win_s1_chipselect                                                (mm_interconnect_0_p2_win_s1_chipselect),                 //                                                              .chipselect
		.p2_win_s1_clken                                                     (mm_interconnect_0_p2_win_s1_clken),                      //                                                              .clken
		.p2_win_s1_debugaccess                                               (mm_interconnect_0_p2_win_s1_debugaccess),                //                                                              .debugaccess
		.start_s1_address                                                    (mm_interconnect_0_start_s1_address),                     //                                                      start_s1.address
		.start_s1_write                                                      (mm_interconnect_0_start_s1_write),                       //                                                              .write
		.start_s1_readdata                                                   (mm_interconnect_0_start_s1_readdata),                    //                                                              .readdata
		.start_s1_writedata                                                  (mm_interconnect_0_start_s1_writedata),                   //                                                              .writedata
		.start_s1_byteenable                                                 (mm_interconnect_0_start_s1_byteenable),                  //                                                              .byteenable
		.start_s1_chipselect                                                 (mm_interconnect_0_start_s1_chipselect),                  //                                                              .chipselect
		.start_s1_clken                                                      (mm_interconnect_0_start_s1_clken),                       //                                                              .clken
		.start_s1_debugaccess                                                (mm_interconnect_0_start_s1_debugaccess),                 //                                                              .debugaccess
		.vga_ball_0_avalon_slave_0_address                                   (mm_interconnect_0_vga_ball_0_avalon_slave_0_address),    //                                     vga_ball_0_avalon_slave_0.address
		.vga_ball_0_avalon_slave_0_write                                     (mm_interconnect_0_vga_ball_0_avalon_slave_0_write),      //                                                              .write
		.vga_ball_0_avalon_slave_0_writedata                                 (mm_interconnect_0_vga_ball_0_avalon_slave_0_writedata),  //                                                              .writedata
		.vga_ball_0_avalon_slave_0_chipselect                                (mm_interconnect_0_vga_ball_0_avalon_slave_0_chipselect)  //                                                              .chipselect
	);

	soc_system_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	soc_system_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_0_h2f_reset_reset),             // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
